//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
G9ttnnSgl0sF2nTFm6uWwqFHiKhBoJhfcKAkaxchzYGbOraxuhbU8ypVNTxQgolu
OaLXdyzCNPlRGtgfLRdp6zpkMWUAsH7mLLkG3QYFB06LgCCh7wM54TJ7f+BAcGYy
L1295bVtTslhutBlUCfdfGkcTdCun6hL34G9PHp8C0J5KHe35Qs8sw==
//pragma protect end_key_block
//pragma protect digest_block
RonrVnQ/ODxeu9rrI31k9DgDJ7Q=
//pragma protect end_digest_block
//pragma protect data_block
B4BfCceadfOZAnta7kpVb6QqLQOicc3mGaDuIypL+KPmA4rcsDSweTuev6BlWAIV
9pmZ1krerALrnVTx+1R2gd2zwjfrGzCW4JC2JeBQNiQEuWsI3KmQnTQuALZpBgha
HnKlDVnkNGe7XBn3hiwlzxr4uA8WA4bxJXlfJxrNeFPFw0owv5RihicOTDDiB91L
eZyaLjWsivAwL7bIl0qkleIo2XmSw6cK1qARNDau901JpQMe7UJwkqDdANlfBCtB
D0lR8KCVAX6qD13b8wNzVn9H0kwtQS6piNqg+CB5jNe7zONClC29jSO2BuwZmMut
Oyf+RPamt+LZVHq4NCScxA==
//pragma protect end_data_block
//pragma protect digest_block
aakJEy3s2RhQf0vjilwIXc2yZx8=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
AvgmD/3MGpz6SK5paLtqSGFiwv1ECxwKxmFa2ojFpIvlTj7XWy/vEqVQYG+QPTVE
Tjjig0xD+ls9pktnZpDJS1NsrVHG2rg01XyHWMEpGs5z8AkIlSQa2DNZL5YCITow
pF94pGyRG4Ug0xkOP+8CSo5MiOnAH7nqtDHcd6MfPokKxA7gdWJYgQ==
//pragma protect end_key_block
//pragma protect digest_block
DcbKornsNkor6wBiuhErxV02ULc=
//pragma protect end_digest_block
//pragma protect data_block
trjsTZBsqZaKKU7qFn6/OpQgF/ao2EzSKeYSfhWe+zmGxRmyJeREzcRyqVSYv/Fm
0lSFMB2ce+LRwHeRmusbwDQ0WH8JAc73/0u3nPgA930sIsegIQCrnWuTJcLEvu71
FbnH4Olaw3lbOfbE6ZQ9IAKrJO3eWgOfpkIeokVve2jMoyJ3vy4FmfTah5irxP2q
MDCZ4zVxfU9wY4V+fBpwSMKm0k/CTAocs66ohUCnd0LJex0zhNaGOReemwhdFMOy
eMwEWnjHfnXLVosnOSilcQm9pdgXLSBVmbffMFQo3MNH99Likq1hZFAy2UjwiLI6
lA0Ekk/VWWjLJ+3lRsYMsw==
//pragma protect end_data_block
//pragma protect digest_block
H5OrBoHAqQVmOHYthQduAkswYH8=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
gRLFMMdgzslwFtgy3VJIh4dE+vzsCthrJA30Uv0nr32FEMc89ze088AQHW0zi7AP
iGRKjhEAVl8XBZjBKAuRPoKbOVwfxg1qhxcV7r46kLMFBlMSoJqYeKk5ymZRNY90
x16ngHc/k4zAuZ46K7/HjrzdjcLJV9rf9icd/16nzQ5YhHKckVt6zQ==
//pragma protect end_key_block
//pragma protect digest_block
MUjBWj2v+itHFHBz7iw0ndqboAw=
//pragma protect end_digest_block
//pragma protect data_block
+Y7h/pl38oxipgKKmWV8Z0HOVclouPwYYi0sAoT40rCleKAhBfiCJNo2nTMbaMU1
xXh1ooq18GOok+G5HvpD7kU7ypV/+7ntJgdXUBPDDY+nwpHYfKKkRfQYoG9yUgWz
wziqCQIIm+6qvC+htoPX98tde/+87DZaMXqqcqey4YndgKcjcx0ylz4t2qIOR0Od
N7BYdUaJYSubXzPYZya6ej2eA1CneNlUxt5zVh38mQZQ2zzqrDs3liNRVAIarG56
gXqAERM7eH4TvwCZw8FgzJEpubU2qiFiSAc1XwCfXmok6cbUhK4RfbdkYwrYGzOE
yDwR4Xic7BvWtIBZhXBXOtwvXNkCxiQK/QRkWm8MZBnvlo5OiFTmhDnZebSpERxX
//qZlMj6Wsc5XowSDnWCTh1T/oPLwmmDnm9D/LdEKSJSw+WJ54TPnSzHkbF0TaLa
y0w3eMtmK+89ue43MtDFlOMUrf4QeSs4rawgLAM9WCdjlnWYfdsyPtSrxefXC89P
izXB0NJewzKqNG2C5Jy9nB/ODmjJS8oxAkoD+peWH3tCO1gjoUKXkL/B1vaTzOda
C4zvWujX3e+lYpK7zuAuBuuWqRs4HcukGEwFa2JXfu2TSXju1g59QucjGB8ENkdy
N+3IiEyt8B7CM01I60MACY5W7osx1iZgUHP0IoDjP1kOEuxPYASBlf9ZYLrAQ+le
ko+DTsRNJwbbS/fYu8ocJjhZbdCkR67nVgwzXM+eeIjn0gYf5OwUJ1W0KOifNOsh
sc0IsZZlRdG17UBNCJ4hldkhwSaynml9YItB0SJsKaSiHpugB3EbgsRroRTsrMQm
fFGP8oH9nefqZho/BVnlcrRkEOEMotOZjHIkRHEUZFG78KlzOYHvdh+0+p+lQ3cA
Pkoo/rHQ8kraDsim55UjHiTvfnVk0jiXtQ+sBCEX29suNN8ArvXi5akuoc56+dco
ehRTczf4BdVSStcje4V2JheulAGr8XbbTJ3YmVR3uteQPN+Qt7Q4iuWQmbb/MqCT
9q/xroY67wJgVEuo3QybFEp61ZO4T9S77OSOzcqDP02m7QcfhYXSJ+zNWy4A6tr6
lQCN+Uq54TaQK8ESp1vPL+mHFqNtXMi4RmyNmBRrqpo2lDf8gUaAONasA3MupiMo
SHyEEXXvPD50uZ3qQnX4zrKdotvZY25oiH8ARvuhX/THaGzmu5b9SdAFA+QYH9PD
GD1Bm5IjqbJ6cyNwpy3/ZnTxJ4kIgfM4xujw7Djz5HTeXY1mGrk329MUzCIh7MYO
1blncHBHknNV+F6mk1NG0o5+IT9THw0gujVztAWsTlPy8RnGStctkN8+XQo4P0NB
lkPpU8PkJkgCzsJwtIuesROok7YDkaG0rMEwwmRd9unDLRx6dQnrmwKAUNwgd5tM
WYsPiEX5hWnXB2nBd73hSEwtCFpPCeU9KG6o5KTmSron4DhGqaUdGIE5IK499Jj5
hbJBty6ZebnRsdjbW9tWiKn6CjgOf6pcR3hCV488JU8Qf6wj/zZKhWcS8e6JCZiW
GlqrHv+eQqHkD0JYCqtaDViq2imqDoh80SU+xXqCqS3iTPfVsnhpeqRh1o0jd8K1
xDdNfUGYmZ/xIwZfbKIP8z5gIKu7WdBaCoCN+FvTGDJPJCnGJemfscZXHPLrxt1w
GrTv6wO23EyXG4Jx3BOQ1drX4nHMUxUMBvDKcJXYkj3u3Ry4xZSSE8OafstOsJmL
XQPV6yGVftQE+z17dgtgxEA6Zc+S87A/YMr8RDWBaOYwm0TjZIYnB7dIfIpjuT4N
ogNYOFWo5vJ9jehJB7o0mKH/TA4UM9r7ROKVl4Tl4oDIuFQ1SBJNShz57CsQwUhx
nhBQUEicqfZtkIPA2qZmBSUlanB2k34FeOCcNlBeYygb6MDnrAfV+i8O3CrZMVuU
YZkWP2jAJVpwDVdsws6F87URS41U+TcgY/SOp7/c8Jr4qH3nBw0kb9doEnGIvf3F
Bm27tBIXGhGc5zaBosHlTgjY9E2NCDJxom/Xg8C7KuCRgW4ft27t8+Sbfa0o3Kb4
hSM86GcRzp7Sz5ZMyczlXFT2rOq0SYvksVeyU6jlBEfjXeK2pGW7+ZxZbG/pkHLf
uBISoF3eyUY/OEYsAudTHENnZp3n5jfnYCGsOp68fLefj55Eyz2FqXo4s2hYSBr+
WI6WSlsglD7Wp6dfUmi3kN3U5nGxNKcw2XpkpEA7jlTQzSRwJTmmL4tbtMRhcgqD
4GeBjewHvvXjvwwJpX0N+bnk6QTIak6g3cDeGqS7j8TDBD0j1jb+pypPhbSCyMWE
OuKbOzXvECdTPc85pZ1ZVvqYsQO19zb/vTq/oezzRp9haDWV/qzLB8HHjAdp/a5Y
HWc5CkpxwbVFxtA+DyYgl6O/NjKwNu4oquuzQDz4LzPuD21Y2Fcf6kvf7pRK9ntO
FQKhqQjjwIsMgSRAzw0GEjw2JPNkku1swEQak1NtB7kc2MbFcagrd0GiFuYUepY0
DBr5NyE57jQlT83qc4pM6ucrwDSe09Pt8d36CFBEqFxtYeZNHoXXNwG0tEV7Q9tv
411ccCDkBSRNwu9TG9aj3YZdRvMKnSqVAgGeKAX0TSLq1ksXG/dk0gqlW1OZNKR2
oRNelzK+0G3cNQ3F3IEoHxRnS1UfnhkX1Z0XhQqVW6qgM83cpQUw6gAHnmjjhT5B
2CNaedIJaT5fMFdZhTgmkQ0OlIk8rnzCHiABxBn83BL2DB3Od0/aqK5L9IBDkEeu
KLUsMFGFuXCrE+Bjp8D8VkwG4OsotIc1oAN+WcE4bk82lH3QhvFOOEiWv5DT3HSn
GZ1EkOML30Wyjkkrzpp+zerRx8WjVdH4B3VE8MTpFZtKpLhX45o30E29EEhwQqQQ
gqHfUGhvCE8Fp1jZB3CNnI0qVyEuJtiNUhqZ8ZNPJd+6JjKJfR9ZDnYDE2Vr173A
lCJTGDq1DgKD/ygiVjVwBmduHSRjzHv0IbS8/nJpzN0Ya0yLKLO1xQwpJt5gDTlD
qmgk4/POO4cxnWkZm5IZWpuauy+i2pSdPW6kHxXFp6Z+wMzbO1eIHnCCci+T0sj4
nZHhDHWlO4QC5pZFQ9Fk/hBxAvC5EVtTEZWh/aec3wfBAiJy3G5ybtguQKkdpouo
WqShlP68F7cDUSwHwCAF0jsJvrwV2POCaL2QuWq28TajQ6BWmPtoIBRj8ORTmXy0
aazhZU4hT07aN8dcNdRjE0rfbTjF81GpOUHJgbehO87KTfajd31Jj4tNitGVRT6u
/P57BLwZlIFy2wkD9VXxwJRGax06IIB1PJUuo5YtynJ3gdCJw5J0pYJpkRx9bmln
l+pGWILnJP1snqorAz6y4k9fUx2vIr85nfU7954Z6NvvISJjzhg2spJuxdfTYoZ7
TmSfh6R4QyDGzwIgFCptKdxKixHvgwU2eMuFmP0yeIjWLn4dHicCnv9pgMvcsSRM
K4ye3JjXargSgFrYcgeeqOoCVqlQSr46egr1YDStaCgZ9MspSRCAT6iHNdZlKqCi
BNrlm1LbRc0Iu7/HFKr2/NI7OW0glFBSmtp9PrxQAFaowH/+HIW+n4UTllt4FODa
hJ4eiyANUxTPNTETdUojwc3V4tumonUvGmUAaMjycyCBnlQkabbofmRpz5tdUUC6
GP89pM7S3ppiRxlD6udbZb8SkzV11WQgSXRsdKIYA34UgG+ll9vYDNqtUDf1eWNL
0tiyWJQh0HSlswFTY8tGXL7SjgkFmI3aZfvzM+G0VpYSobWrcUG8shC0R33j31bo
UulnhhdU9TRTMpyXQAPwEX3WTqV770KykRJ3SnGJHl02d+6hN6o9Bfa0C7bA7EKG
yzycIONtNX3Al8Z2QqyhdTBEJ4/MnZ6lGddEH8zuYY0C/szFDbQaJElHmygJjmxa
ZeOVJfV4jiVguqvbcP9XYQOQBx9QJaXTdlRTWNe+pg1SJmp4xk41j8raWf5mHL3O
TK6i8INubZrhx6cHMiujGcuX+wKKRFY/Gvft13Qy3ZrMGOpj1IkL3yYwE5Cme5AT
V4dY/gxhcxme95ZROLp/ItRE6ID3/f2SsySUx1KQOCMFGzhb3i52BB+oFv1u4UAH
xZPyiVqZZNfRJ21nAawSY0BRo9IiO0Dw/+79afBvHFLLQzRG9OvpmGMgQ3f0/Q5/
1eDXOLRALLbzxd/iMtBT9M6uM2bgiFgl6SfHaM3odxVvnvbEdhF47bOUKRM9WoqI
czh+KRF9kaWiabPMVLA0hgxH+uwcWrQDa1BR8LMzNzhPOtwzK8Wh4hwV5Cu20/7v
ezAW7zvd6g9dvSX48m+BkewNcXDcQkm+jp/hr0Wi21Wlu6mxDb3kdDFXe12fSupj
UfOGJ7PzJyqeiSyub/mlpgFcOSWAWFNe839MMvKCi3mdWhjLv6rCoeYCE4ZZhS5J
JiZefWGcYT93ELGKJ64NJODKnnN/MpZQhIbaXzi8H+2QDvs1GcvAUKAcZVgHNxIN
e5ZtQSWA4sP8h7HcqtKFSnAMBOD7AKDKIrA4DdYj1tWQc2VpZf0Cx5R6YvxUJZmT
u3G8ud4oFg1sWTcsZm0051Aj7gT1Y0uwwmyKf0eZcdQILY26BsPd0o4aYAum6U1/
JplRl2c9VCIqMhnyAj7ST5aFcyfQL0ROiCpIJtt78wol+tZQSvktpgvwzxPwtMai
UaHt2sZjl4DXec7X6MOJDi+tbqPqSWkeL4if35cE0V0MzMFnn0PCFz6VFmwzqiey
c+7sbd1vkkddcaxgk3/0eAcUNB9PFWH26jJ8eMKYgwyCV+vDazJCHs9TVD8miqEs
vYOI60yddD/OpqDgLExG6ruvQrJwcvQMWDRmdOcbuUSLYow1shicSjR0mYrUMO9f
94lTaxpJTWf6RQJgAj3PROf7ALvttjTtkvtWb9Gsdv29xXJuYF6wW/AU5Zy4w2pO
aK2Hf+ZtmHj76DQqV3JdPOuFa5QGlK+hCHFftJILE90Y5VVuBrIV+nayDPA/nowl
Nsm7zuR3SlOrgInXPbNYUG9P0YkEpeAxTxE/xk56OXHMYA1ZoQoYakikxlnDdOp+
vXjZ+QNklWH/qWoZ1025WjIKUY6rei4bORlL8/48etgZGg2XnPLO0z1cMUd8cpOM
eGRwYIJsPGvyL4tVhev3nMxLpMSg1bZ+/kR1T3jJQO5DaFdgM9y8AfJ8fxLyjOzv
nydCzGHuKzYKzq6k9vy3chEhO1biB7+dpc1AYC0unJBNkX6X6gngcRYAwEuU0qdn
5UYZTBc1K/H1HQq012QKdw5fWj1k8rXE0gUocnbDT/IjH9fdJNxlbdTcfUUTV7N9
FzlCoBLqE4P2AABlANCgJ1qCqWxDJnlFJSqXLX98EScqdHcaYO4Cnhi+Xnx+ryt6
uOuZwS5bBbRw7HYf1VIDs/h7nvLctpHs7L6uH8JiXHMrr7+UY7YfPdQJzn/j9C6K
TuMgRDUxAcyZal/xBzN/iiHZehhWtNSvPhhO88iaKU4mc+ZH1A/pA5N4PbI1uuPM
JqzcUS9mEp+ShqsOaTxJWleXgNVbvqPyKYUjHb4jWwutMYaTi6I5j+HuYtR1+cd7
OzlkIbJjcD4oU/XajQXowiaJwF6uB+aHBILhGi9J/tXB8JytZ8wmR5HGJs67zZf9
e8U7BlgUj23+qEFKCs38YfcXsUOLk/csS/N7Gq4+VfL3i64I6ENT2JAh5bE/RWHH
aviyYv1eT1jxy8s9qALeF+FjSFKCw6hlvyyYhO7RdrrMWHYyO0SNynXM1SbjG7Oe
5ECcFu6xm4lWGsoMFjjd2UQihIk2qD8flSiiB2WpeQB3u7cHqbTSSsK/VPAEEv03
k6+c1GWLE6C07joIds+7RjxbqY8AZHteeCPL84qpJM7xTXQa83eqJaSThUgfA6Jp
pmVSeDx+nPlAGh0JLiugPSZY76OreLeGOp1ZFNH4is5agLEvvxSOqE80wNBxRPqV
tOnQ3TgCv//pJF48t83dhYC2c/XSJGqOGpriXE/w4/59BPsJ9H1vxwIdZ8Wp195a
bi/eSyFUkAgX2zezJPc1efyhe/o+iazZPIkdZCTWekz9N585RnuAUBrO/iVYIx0V
qf54RFO11lP0G/BkQafbm62IEQsStDyauXfmPj48TKaZKLCvjLBUNDqfppyi6pcT
KoyaW1VHJvLcuGGwLMAEfrrmYiFt7RZ7XW/+AyBThAi0emRXLnj5DLDrDYLG5TW+
R4V+2Es9ahVXyg0bR0GjKUcbOhrBw+8+yuZeLFZGFityINRnA+qyRnQ755B6nCKf
hBhnIWb6Y1dPlwdd1Ne/kOjuGsUOGt3V0Rq72G5nvYJwftu+cI3y3bLSmZCD1qhF
zBBTfOaZJyjOxUGFD/xkt5r6LzML8S8TyFY/5kJq14kq7i+esROyjKddo9RAPlqj
lUrmdk9n9DN6C8czP05mekZXNMZzdBpllWdVOpRESC4twlajb6X0UI/lsoKNFjzY
7cmKX4+RA5dviphIJTuA4PdRUSaGMgkaToWSOz3o+DRDWSHRmUNa2wJHRCdmTKlS
3Y9LtLJEnIw+Tx2HvxLXo2GKQUTZ8u1hC+dZihhjSmjPGaSuDt3G9PwF2+NTpNmy
BB2h5IwDzrogEmSjMLvk7KM3PkzGZNSIionhWL/YmhgJDjTXz/9z4T/EZ0UO7Cp4
elqDQTYVbqKajAeN24pw3PfhhYY+4UFRXQDEz10d0v0nYCEk7UXrQ7jPAAWqGh7t
c4iRa6ObvmUHyecxp1fLcAuXIOD6fvjmYTeivE90pGpYZ0CaF4TgJHZhddEyjGsC
sPOI25CcihxsCgRhUN8FqKNsOTJDVkEqlqIuTFeckszGZuQJBpF3UiW3xnCr0RJ4
ecuJEpK2dhk0e1Q7cuKLw4t9Q1mcAa0UeXUeI+OUbqtey7RGr02jT6tGnHHq4ZN0
O9nU2mRMNXKzcf4zhp57Q7gbR3j1fyblB0ZO8vJPXoyhqQauFUY+N9KR8dPXEUg+
2K2hknnnSv6qY+CKFeBpo/1ODxNKhf4g8MlcdZ9EEUZce+vxXh935uBe5BGkUr7S
DoF4zKV+roaCmj9p4KudwZ88xuFVDXBbUf0VkxnsbL1lMu8mg8b2U5bwp0JBb7co
Mbck8RQNbClT9OkvICbJsibxXm3QSy9dwZn3U/O6pwHJ59b0WbGZP+zzdpRJITzk
LD9l/ICAd0M+M9MMnVmkGhv1z78URZFbV/DNKwccDyQsyh+Erlof/P9hUkP4KcWS
L9p7o+1kALDnfBl8Trh/dqTUBWWJrupEr1aB10P1kvr9HX1dFAxz0mz7a/YzWWbp
XidmbA8klixFXGnuM+6kCFDtiT9qOEfds3eRgInBQVsYQRe82z2QVsjfoj7R8hgR
8VjdxiBN73S3EzYpHWW2vKWgv3OfUuXkR1tVZF7AWJ5XitOZe5r30r9N0sYVxMl5
tGUVYfwEGARsMa1NpGfOnSyCQnWMQaQ+gwoMdDoEZZC5HaQD4QuhuXEyRyrlC6+z
WfbpJyJh2axyIKC2XxjdVhalYdixJfiPvjpWWzUZwdH8+/Z8TTqOgl8eL66rdZHP
RFMQ0ksAiktYCo/SQoLQdCAgCNtC0y8l0Iv5Oes5i+vvf96LCV2WIIwDdfvEIIAF
D7bjGZL/EjI7LHfwL92G10oyZNxoL+Xr2B3nvXeKMWqGgcXfBDiAM2qadmrHcZr6
ERaVsNyDG4Hxv8oIIIjqBZScjHYbI9qelSZX5G2psjfqBGFGTwv9HRW4cDfcC8Ni
ytxzMafuhkPlWG01SOw1BTkKSIh256Gob6Z6fmIcPLQoi93axqtnBKk4yoq48mV/
B6CXe89KavPOsP0CmoMg/BD8uACBE+ds7XMNJOjdy4VJrTSyftgjduohl4uAQgj1
JKhA2Hpe0lGNpU5xb9fe1WYC/krReVX7jPjfNblNBpmWHjZdQ3ZoDvjWNcGJsMJj
ZKMzectZu4dJdzU310BJZocEfRs5F768A4OKZkMNe9o64Zj6hid8Jdw/vLr0OCjF
QxnbhNi70xSfRb/njv/IkTC+iWVBvkUc2rPJaxZQVrBrwCuVHtqZAlRtuNbmMqOw
BlN/vKJ8gZvIxNYU5Dfo895LtkiELKACvBd8xrfBnNaLUTHBdqtn1I0ker1rOrOx
W6EFS98UJCaolQe9JNose+8FwvFWKjNEMOTS3MFaOej4N2vmyvzQwAO3KE706SE5
OdS6UZTrIxPDTCmfFlsMHgMaZoI4cLycItVBCuRBnfp/mLLb6Fir/GdfE4fR1vNA
Ear67AoQ81rwp7vrCnq/mldB+M3XahgRqGfYhiAZo0tsPtoss90JPDa9uIZVJfyH
p+DdgLjtmOh8DuE+BtZGjqp1Hl8DSfHfyGF8pJDl6AUbORPuNhSec4FdgR688LMw
A9q/i8OyEwqUVl5TsSYSOzOpfB17rN0EZP0qDZl9VnpsxotgzvrjPKlBMMyO5BoJ
pEnl9xFt8P0tJWsOhg8y6M2nRdnhm6OTnF8yVVY3o1VlhasxJK8cowAqBX5ZULia
OgS0OoBWIm65EiXNCy0PfDF40B9cGckak4VXSlN8Yz2yEytplGB0HMLS9hkXGJik
XBXuUqoeQCy2YOc2P7hJIwBx8+Q73Pg66DZrQpY1vxoK76UcK1TLwuI1vqrH2LTa
PQv7r4kgdGtmiV8ONl1O14ylXmsuOYFJI7xMmnQ75b0tAfjTmKUrSfRUJGjiaVth
vACRkUYwWWc/wbAfy4feSm7yUH+EePgdbnMiUiU+wFAj00bhHTndqhypSDCTgor7
ZrxBC+BAPivN/o5YGyAQk0dpFKXjUOmWLcY5vP+4dgEbIKnHi0PDyzaVcUWAzZth
lyOM+BaAwv4dmT9klJIVc9dLAba2LCFVLyimkvE2s+HPc08A27/jP91drgft0OP5
cQcYbOWS1OJ59ELRaTZ/wrACQ5x+OiEixXgjfXSnBxpi8kwnznEiqPd0uuA/xjjN
Vu0S5/+sdauoLr/UsTeaJc10PHJALREyH5UhtmRYuVZSG2H1hLKlO6UqGV53zf1i
JkKbzLHIli3QKedQF1xaaIIH/nGau7oaVdRljTzoOsdNubx6L/tlcM7rxToSTWot
UfNfYS2UakmbUcjM2cwI5RLEkD2N/jmreb6OhtKX/BW50Hgl4tWDj97F9fcLlDmy
qKP0/YrRwSZGE/sHlGSKAWPnewhHe+H20FaLwAPKdZ+P3eUgkwaGHJ1lMWi6jeH0
07v5ILkfDPuZBUrMJpPaN/D3etkHaiX66zaZCLJ0fzvcxvwwkLHmy2CUSCA9OftX
buKCHIlgXK1SZ6oAivb2Sg4Wp7/NamJgKg3ZoL2JwAc38h4H7lLbJG28r6AxPesM
yhidBmbLdeMzt1fY8iYFrc2op7G2R5wMLFlxjfTbNNlklgeZkxnRmwd2kvu1UCRU
QVnMgrk/X/REPV+UT/X5nBn3Ic5JDfftOFOAqOH23nPhe2HCRowedGkcPNzb5wEb
aSZyTMHV+bBgENg4WLEXrZVsFNW+e9UaIH51dWupmW60p23lYOKBlNrwH6RHCdCJ
zmPH4vJqdKaOIBOrc9R1UXniRTgRjaFJnjiclu8iLhtu9AZAVvy8UnfaOZrC3X65
yOYQuWFyNNxyStC8J3F/lyS2BiHUT8pDANeQalqIfXLPUeYRMQcSwuEtDOTcbPXI
IhyFVp0uutyprM9VJw2TPDjEKNNUcViNSFKtnM49pOUnvMDd4MZJekjO1Ko8v3UG
MYyya42lcnuAocefx2xTIcst5W9oco6PaTVLJ+HCxd39KjH0HTN8KQjiHVms345c
afpK+xpzUUZLE41km4wrxyh1dCCVrvJDMgAlgyQv7ICtWWYEuwosl5vuoOPuPgP7
RMRNrsylMGkaplF+o86tFN2yut6o+in2pSbS8gZKWj1x1ZF+ogWxNFi7O8VcLQZd
ywj/0yMMMM+tcUc0JNVLj87hGwRwQIIuvyRBgOdYONeeYaJPnjuuLW6KHas2q+6T
4Cd1ApQ8elmQdhpNjkB1gbz7WkKHkMfizophEr3MYeO5r/DtoRyFIccOAk0i7wSy
2D0OXnfwparcPw4ZQytsAb8ofqibmwsLYuVEvnZTc/XE5YKhao5iJro264zWlHSt
nZ6UlFubj9PxBEc0HgIUOsqyDSXksYpIzr17xijlgkduAEcBhM+U/12HAYi9Qwf6
SG/Q+MsY0qbPmP//dNm0r8kRcycjC5QSJmUVNK4ODkDvs3GCZTni3fXx7VYSDe0S
UMGkBegxrsMB6wkluScXNTKj2Af5J2ql3NjfWjdTA6mz37ZrB8cpkZFwAob76OEC
i7fSLtXgVsnu4ZBRj3T9/+Ksn1f8hGVsRitldTAkaQuDIFUjaUpucoZkuEw5SBo7
9BtIl7lRF3776ZqzuvcEd3WyYg+oIsXyp2W5+B6bhVTPJXQj1EnlL1mexHOYXgqG
o8qTfWtXIZiK2q4eM00UZCfH5TOzR/ernRDBjChexNQpDiszdaQB5tJob8aAdMpR
M7fSp9iPXB6dUvfhRGIbfg9EQIHSrAa9api5wov1PwKRn+cYggzE6FkSvrB4ZQ4l
kuAEbuX6aUMPEy9hN/r7AsGMLFcnlkVJ2Nrh6qzX/XIcO0xoc2SJtUItYXw7KKln
+/8MDaSn5QOkFyMRvzNo/Ewjnkvcn3TTCsGLtxnVs/9vCxlTVdLwlG48ye0qqqi1
xg5ez3lCWRYRbyJleJtr9LoOnrAiQzQf0dJ8lg9+XiOriZSjXBdW6rIFBXksjM42
PozlTbtBbS8QvXCmJaWbX5E8ynAUK23ESM+NT4mzXOFI5F0401ucBBOx5WaSDmg5
mZ31YVlpq3a60BP0GKMYQQheGnoEaDZb+pTjCCu+V9IS1U9TUSuwVkLK5iQenlwN
swYcBtKL7kz7m59HvrRDzD4+7KlSJ3vEJNanuG/6zhi/XqM7cAkzo7MfFDmcd3gF
4moA0tksL3IRQN9OZ7lyFBQJpAJCLREiNtdM1dygBnrR3/9Qrb32t4WiCJVVWu2K
E//6dEgn7Sso2odlEh5YMyNyR+srhKsH1EkDvcJQOSPvyPTB44MjsT80dFk5wLcb
ZrA/q3a3zS8sZhiL7y1ZPiDRElAlJ/HzJwx2gPo4+BoZ4C+mbw2aKNZ4dPmuyq/W
oYtowwEhU9xd45/6uvIYk7LY6sMKWw8q1QrWDxLI98WkdQqi4H5kM4mHNcgRj6i9
9jG42yz5gD4Vu2WIJZCnK4IeXBPOOpoiCz3fCl8Xqpg/j2UAsPd1UdROpP3ZPpMO
xZKJDQF/CcOdf8fBKZGGIb0zi1b4Yi7S5SOoqEY5mESVZxh0VURrbMAbwa+Zu1QI
kEu0mSnE+c4bLnxKtDWpDOOqjhN9IaX15wjM6eJg9yT41s9aob6naYNMB1XEc25K
i145Hvfiwo6sv6/cTdHL9KSrbp5yTJVByxKHAYskg6WFtp3+JjCI7eF1K5TpfFun
WHzeJlHZmvnaRdgWgVunoCiCxpoNIRO6YHR31NxShS1QC0F/EaYm+dJPgqNZ0q6Y
WYFfUU60ZaMuvYSn9jf1JRdsv1t3Jo4q1lkI5lywieBbxG9xg5xT4j5mdgJkfjAr
GJo5NU04OAPJQhGM1+qegVMTmaChki/ULQ1xV137fAxOsKZz3kRStNOlIkFdOlFZ
HqOQxfz1QiMmqAmvm1ruvO66CpKPovFmKz3UYwS1c/oDFRqaji9Ykf/p3dnwCh0j
To5saZTbafynqr51JdtglyCrzB9Dw3UpxzRUnc+tBy73NKaYgKU/TfkMmT80SEKs
uNYCcVviUW0Se2D+1eVLpAT9mrlbN2DgrANcRf0TV3m5e0xvzZ5kYzz/Fe5hh+YR
ESutTa9Z6q7jGj+JEy+IjtMSKREaS73IwE/1Ql73BBRcDzMYLZDcEXDFCTo65VI6
IyIDJ7Ca60RHQKkErsjzjLl12+sdQ9gOaPYqNdRP0lnegnuzXRjEn4aRUJfCOEwY
Q+rR75u5lQDYadojTOHTcTqmxGkfrTrpABib9zVx1tpDVunv2tDI1SxXW1YSUhFF
3Wl2kw4jW5kMzEuhqzNHpwEm/YNej0jSD/QCvbg3/0JInmhLrfWAMGwf9TXzk8PS
9aT50S4h4b3JGYuhSajFP6FpRliGIYYkp9gCfyGW9kpNrZaJcqGFupMcYZObymYZ
FysBH8Koi5+4B2kt5GQCptSmENU5I3wse5oSg1EUMKTuFFblHsD6fSjY0QPU0Jqy
TbHhWNvrab6LpDcfZLgTW1qi06mDPXRVWLkOgSspkgfcDkQEeC3gokBbfOjcJ6/e
sQDeo+xl3VmrBryFLDmL1vW8Yj9y6S94hIPfhLPE/1DC9iL9L6Nr0XyB1TFBtRqP
j1juvTuk4FyaQ6MTLWF/i8nXu7axMoCE5K9joEZIbWtEsgu60l378MabLT9o8Ve5
wZWkPbznDLuFKKIsrxqL60XwRCUElYQ7Zhp7HuztJIuH+P99T5xhwSp02Ft4pU5y
22c3OJnd0JJK2vFfLx4GnXYMqDVWhhekT06MKc+J2d7dZtnQ5wjExuoCMW9o9T8n
ssa6lxNoRDZBXqbZFA/w0nFY4QIAJlPiaAMrc3uLTqIkDejO/fcrlzIbs2HeeVaZ
aPSMq8hGR7Y2rR+2m8pFXFDknzVdpZtxBME7XNVTrCO6CdaEvCmQpvxH2vp4Y5er
FxXIZSHsR9VAJJGU97d2bNKDfiTcIVt41M8P/B4ILFsRNsJpvLM5ep7EHxvDVMmx
9RWmBBWWRv5K9APR2sYrkrUgZ1gdE3/0KZDkD0YViTSUZrNNn0Jd3z4doobBjeNy
mkVJqDKJ1UQQ3j9PAK79tXyIpzl4uTsGUdU+R2nNPT5bBvL2Csz4cd1LMMAomuJB
zSksXh0UJNFUGHR4sSrbB9jGb7ijrLqHZBncK4e6GSnL/aCoDrobfDzodxeMmVRf
xCoYij+lZUvXwNxuSa71BMVvt9FWZDVNyEWkzWr14xtTSqtBy1PCRSyDiRBoawXB
aF+LEWTAjXoyApZdlNDTDS0x8PYD19KIX7r1/qhDGsDY+i9mpz1aSD+dXEdDmzg3
txLi3VT0AJApAWhdEQd552IxMcyFBrgJBuxD3fhselCiSMas3Ft17kb0+LCi5QiZ
0sfYmc7/8g6KnuNnMeQey0nbqNlY81Bytx9QwQ52WL4fBmqmqTZQgPx3d1wwRusD
0mKm2Je5ZyTkuOuvLjJU9kpKWChAT1vjk6UndRs81e6y0ad2O0/nWxCOXnRCJmIl
tOdNlW/8EXGec1S+O+/4Geo2dFJlFYrnDUjOmajXTv5Y11p7Xk8pZSRM5BaJUYrh
qGTaNcOqlUDxhUBvCpy1x4zPjuJGKC+r2TIK9s+PUwfUT9hgGmzxTzr0oSZElhUs
Oo8nvpqAH9DSumF8Ga2M9PXDXHKge4s7TpN5N/+xXHn+WpczB9lu8N618OaktUw4
WMVTrw4di+yn8YAsXYP6xgBsQ078ZvNqBj2sEdEspN5BOM2hdQablSaEED0IP4pt
4KMuXProvAKaIUAc924S1V6ohxMGk/ux0TODoJ6ZTuoq6+BsJvt5FLP99KrW+wyp
IzUII+BbET2S7ZUpfmw9fszi4Wx8fP3MDXq0gP4vGxfm4uKeSP110DS9TGzT6s6L
2xCoo7zAHEZEU0SD+rlo4DF57AtfqkJuW3J+bQKt5qccWvSTh2/JUU2JFZkpR3VJ
LC6qIBKhw9gRjgAD2SpguS6n+p6zRZAWCFdbVY31aE/K++czrZJFhfLmp9TmwHPj
n1e96DX1+DK4DVWtpMlS1q4HOEeZod3o37eSYJL1vcVC6nXtCp1apqWeSECtDpJQ
BEt+a5i4oOuPN60O+UuCU+r9w67YKlc3XXkklVm7n/VMjZFqpg7jLP5BHTLMrFNi
Xz4+2YSx+8zi174muN9ZBRl9Gcld1UkdpHV03g/01FbC17BVfsK46acDx2Z7U2rL
JKzKd+onus8I3MKRcf3LCJTaqEUGphiAvB3A26/aGdQGrgWPeXRhl9eKYrYHwmi9
BplSzmZWJwGdT0c9O0Dt23sLGWk/EN8TGcQIKCYM2dlw63B90zeu0yvzlnoWoAnh
N3mnZEQXh9TL+fI6FMKlCaqxOESTl/aJ3wrBctZoIQYXtHyLsf50kzKyzwWT3p4q
6GaK/IIvVUgT6k+Sx87qMs8JS3v2P1d6If+zIubG2qGNddjJYDqWkBFGk5d7MHK6
0E/P+YVye+blShwmW4e9OKHjXmmCAwaI9l0iBLjhvcloVKY/rlAQoEyY+7VaVyvB
SBpxQuA7y8qzakN47BKzGj/leiiTEPOvGS/6XemSoT0gZM/gFm0T870mPrzl2rmr
4SOegF2FkXx2fICy8yj11RJfylaOoILeOxyjIS4kviS/4IaO1tdO19VD0rl+iRYK
bWsJBWR48UZr18HVCRIwo91fm0GtEe8jjwzRF1CrZnU2FWbPMGYqnjB17dvfr+F/
6IxOW+o4UgF3cvZ2S1Vj8ACjxqzoOa2JF9hKXMtS9YbQLZSIwOEpqijiC0yFxpBT
GvJbnxlj/mIQE5rLSGtsH5WdArv3Dwc+i736Q3BcGcVK/75fNrzyXHYcu34phb6V
Z6MAFqWW1jbo9ZwuCdPHjRsq2lIyXEqJ9Z5V+oCVMqXci0ZmVyjznfWreJ6v82e0
5R0+yHqbxwFLNjmULGKS9S5hZ0nNJrrSoVYWebbT52s44L8dm4x4q3j4hgSXpgCt
GAcvZ5h1UfngzKcOn0cbakdBlQEGfkYBa+XxujHaVmqN6TF6PEV0XwVIFdB9RDTF
XoS8TMcYljzCiajESQvcPjWklWXazYH0d+mLhbClx1jkQ+IvhQrLR6RVguU8hDNN
dZpCA5x5+vMKJW166NJqQjPFPat78q9FvRbAxdXiWpBG5tYW3eidhcKKGr8rwbfL
mh+l+ckZJSIVBsbKzUQZF99CvKRnWuPpgRXB1QqOGLBrJWi0RTLQvFJJQJHVfpqy
juCh3UWrupXRbDHbvG9vZDp+YOf/6XWG6+8MQSR4iCX8OXkeQMRW4AAZZFKlvngd
tf8Df0F8HW7tIpJrdKk9yw4r/Qd1HCD6LYFi1Jy8OEasAWtknTbdfSwIK7mCytJx
nLXxQYvGScr6XjUBXCWQOKLmektLjq2VsvQ60m/RnP2ltMoINEfBsT3Dw9AWLhLB
4OQmWvOYWV37EHDNQUQ8Eoxs8zw/HDlPeEnhaHeCa9tmwAY5oiPMVSesVE+Vqitn
7hrfoxcCI9dXQtnkffngja8TlotkFOzDYypdYR76nIu5v6murng9shDGSwW8NPyH
NppLtwWZe0nSzm9st/S/FgFtJOOvh7DDwdCgc0k3h0stM+5DAN5PDAeb+Xo41qOs
cFa3MA/0+gx+qipAcZliM9Hovl+x7wcpSlSVXmLDV8I/ta4PxKbsYNUTe8eUiXnI
KclNN7q2JThYK2T7oCIcLC8Md3GNDNkbH6m8UnDvaVSaAgWwSSVeGUz1Hd11BsmY
KGYRRb8tgfdhJr2zpxA1aaN+Uy+gR8H7HDjIe8EZPN7808+D7pPfr/IxAVIRvtHt
NLRBFDN8PMdbmFqTTSgA/XUkI+LHvd68BzroCf/yxI1mht0F/KTpVgFAJJZoJGh+
yx/M+cqmQEjujCDblFzxElmSahw/cwNZoKZ+EF7Iwn5EWpYNYnzyiTHzKgNmWf4z
BPTPQe08pt0lqwHFmTP4Pj7Xqh8c8HQxpU53sJsMohOT5bGv2UV+e1+M5rlZbVwq
K+M/6pzcv2dkhEY1ev7AAUdOT5yR3AXgITJt9Te183DOoxXWVfjdvIWU3uBIxs1r
VoHAMZ/NnK3SySk19gq0Yo1Xcl+8+/laO6gCzR7ODLSAxkhSfSd3FXik4HZgBb4W
fwWjccXdGVJfjuJzMxs63ioxkyhAfwUGXF3t96XgaoEakkXy5+LbTf1J231Sqn+z
WhUykTbDcYzTUN8amOvqrGLS3fJkkOgVKCcVbYIXNvk/+PiFlPaMaZmLAkKXucR1
kORwBaCIAdcPDe50KpCKxpKBadcQneQgfaLifDEjmR3IjunYDSHMFoNxU9vbgD8d
EhxZ0nsxD9YEjyPlIbArxSva49NLPdblWNN1biR/hJQOcolAlA3QC1XVyQm9GFpA
3JWVkf2xALDBojy/oZzREAEJvJxLiV888KPqlqcDS7szZCGqw/fjhaUbTGVOva8S
SnBI94e32JNEk1KOq0hfWZggdu+H/4fgZDWop8Coi7DEFoOFq+bqXwucBMSBJYX7
1VD9byX5mnuD12lHRWhtIFjkbWLFgqIwARDuBCSJgnDhF/JuREdf1C6YIyfXtCMP
R1bqvhzzouaMSQpPND8DUoQsK9547XDNtw0nJ/SBkaVQLSp6EIEK5jyLgkNUbepg
oUcHIdOEoM70bJLFShQ3CtjdOZLcbzvoBTf54iywqz5fyUFm53WJ78BlqurdaSko
uEFrNltiJ6mog8QHsi1sMP+LUvo23RkYSN4n1DGaRfBLgMZlITNO/UFtFlALFff0
YoHq0WfTsQy2ax/8Xx1WL/Aa+X6EVDvPtsj/K3PdFhAOnAMv/VuICqOOWIFW5ZFy
SFSr11YqPvw8tl5S5dK1jnelz52jAAz/8TrlVJ0IvjX2Zxt2yOz9Khi+AGAAr/kP
DIJmqrTjAqm2RsUO57yG8JMTP77z+SKxKJLXqKwK/r8o2oDOWJHuehAMogaBhlfp
EJmJ0LH4D1wPB+a5uzrifWbbkJY/bFP1bKLWEW+hOXEmnKix03iCTHhVDj2WXasl
9xbWPZ9rG4j/IXXzT1tEcSop5QWM6yzEVp9bJ2WU5dTGCdoKGoOTnydLrMDFgEVb
bEh7xy7J8QDOKnIeuIYIpAOKgRdnZwmHC99Z/6CK0HcirwWXn3VHVs73etPuNfbS
M40IrLpNt1AD1BZ9IBfKg3cTd/ZSvxqhEDtBMvrLnvx1DrKr/szGL4wLoM46xNr/
vdNAMdiy4DBVEQB/ntE+3y573eF6gGTAuimuSbcku8gzbPcSSEH9x1Rp7YoVRy4E
7uRKD6NdUyeFH2YEaXgXGiYUzLUC/rqtbjQhrjH+Xbx+vxZ7fTyvGTU3u2C+lFH0
oQQ+VuhKrclzVWQDWsv264btKZ006OAg8Cm2n2dfea+fET4rqymqt6hUCFDpKGl4
OMUd7nDwNFQy22TAJ6w4LKhkFlC1tZow6suAAZ1Aa7vpPaSOl2VcOC3v2bGOeqd1
SfqvAupPbZqcc8POCEkPfFMOSgCEujIOMa5lsr2g/B0616dSM9+Aan9uPRX+Xc96
COVz54cwwSNupTAAGTw9C5HvwXlyHHVmcfIXG+LCY77YmbMLaNc9UdD7UH6MKyCH
+1wHGgmPOhKvQ6Mqyq3Q2xIsBTrmiRIFsrO8Eq8eD04CzbuE3iycRwbLjQElr7q1
GCZHqnnbIk9EThm1x60E9ti4IJVcr2YJWAKMR7Wo0GwcLwI15l3EmPGcbLwtXpGA
3Bd6xDYnu40Y9VB6b8rhFJ7Ivy8LMXzK6exjFeOWAwlqGwH+LuU02DZrwqUg4IZ8
dFKOStUSAFvLsCriS1DOFQUwhi4tg2IqflEobOURUTtQZ3ePueTrbdtGQZBSDbBd
f2KRDBj7H/bg9mRq3o29TWa/JVvinE4nzNGlhOcG8vxKLwTH1W29FqV5ng+eNvxV
ulqKqTd63kQ1HaRHMb75g+dM2EmB17066dP8KCCgflk8F86NYWhKjdILLIge4dTT
Jfo+MENe57pPSwqdVLIKzOjd6p2TyEBRH6JdYZh83qMGMulDzp+xIBEc7Hk6TSzh
wEalzAXvWcWt08+w65wgJZYZUqcfLQGg9G7SPXjL4CkNhpwzWBSwwwnIyex6KJLM
WLtoSV31fWHpWSUbvGl06GLthVn7w4s5TFA7ASK2kI+0m8B8CditOuYvvAIMe7Zj
3axoasYJtpiIqNddXgf+TAZNRGvfCIpeEXkf4xd18CJBvih5zgC11NJIaiypJ1Bn
5sP0BO8Arhh9a6KgWhxeC6jjSENOpSM9Reai9eJO1f+PxNlsOQAfVN66AeabgD2F
lkUUJTQujtRXvvFV9hYSGJkSHx88b3DrDlQ3tdLgju14BZvp0FqbhCeq5Yl6jZ4M
qJC3QFoctrBGcaEdCuA1q/y9X73oW9qASayxVf/R+Ifs5AsYksHzbum+Ymb7nZDd
O2s426nZ2ylMzgDUhvB0SRWA+hageFvgSSCJsJkZPG7D7bo+8QjTGa/5hPKOWqoY
4kz41ticq0m8lbn1Dw/ZFceA8byEekyGMBlna8tcXS2Um3y+1fps3aXg3vPdHcRM
aAu3iOmaSUMtbvG8uXasWPLwQFxWaq7I1LRtaPZ21gAQiFSUYc5178jpj5zk16p+
hThP+DonTyomldioeppa9siIqD5Yigj3Gn8lKuCwVmR/q2YgEjhXMSLVcZlacTpH
rF8uMMa4I94x2F35qp2zyRIYmQ8FovS/z6GE9tqclYDUFjYuD9tjQPPwP6hckNZV
QeU+zcLfX0HWRT8eO+rw3JjCtrblAY8a2CtdwqgR6LNqmZdrcwUob0BHA5Z+epWe
sK3b2DvxAZbajXhdcguqFparHhTbY+6K/p121YQ+Vmu4koGCy4Z3yrKDoxqMWXPf
X8SuoGAf4VYY5g/rTJWgV2pTRP87dYqi3mg+3B06sp8QWe8m4mYkBQAZieAdRqpC
2DIjneDUvR5Y2G7zcfkk4rzL6U6rWoSjKifZdXXG9+zcL6Bg/eKXdouBPTGz2JFk
xAbaKXCGRwiLFrZ8uRmmrJQ8uu85ILur1dRa/CaIK2JA2StLZ8Fpuvnd+XUfMuS1
2TxH20xjaQzG/Vx3lE+x9x48iO701qxOZ8XH/ntBiIEzvy8k2Cm7CImYg7Y/DQfw
2XhWonEKl9jqTrrRaoZGSFaZDIB1bJ5iyw89rVFEW6ou4DTP4X7oS+6wng74uP0B
OUCyKlABz3tviHqK0RuclqBiyxM7Tac2butjlYTj7WbydBnobLTAHlLi8sP0+Gdn
4aCP/IgCOQuSgJZTIw12pRZb70EUSBkhGSS9IV4iyMTm0WlkZ+xKNyIGOY2DNkFf
jbJUB7ZSXqy3gLENQewhlw5a2bJMhGuweb9McRYiBAwcGCwQqGP8f9PCxP8qT1pB
8AH2LYY2Kg8CIvD3FNr2eMgMI3mOBG9ATkCifuSINT6OhyMlult0LxPMGz3JXrGw
tv/TKEA6ayQUYIoCddqAIPVTwV4G9Vhb2BadHDuKBl772ubL250uHFU4c6fpAJh5
kvVD5a3BVptdgWXZRwAXtl6EZa0Tz+pa5SGesyOkus0McJeXmofzkYZQ/KgS27n3
SBiAzhVc6/mPVPEc4NjJpp3A4uMPTyT9fc2HSdeenzNtFsC8Y9A9jgGxUyZsnLL3
bfWRtJk4m46AX557JvTy29u3A3E7Q/adM7QC3W8LJBNB6NoBjiLRnISM1FfKyVZG
sdNKVtYet2RQbmCX2u1afg2AU52XXhlauATrzAnuBuKBe5nGesIMVqbTC+wK+C0+
b46GjcDJ7HfhyRg+EYLszzseYaZc708C25QzZb2a7fYULoZ8quKKEwip3Pxnc/0j
ArDIFEDDvAF/wDpWFqJzRkwsuUBwTJF52POPkkNknSgzaBMt01RqJFzNNLDwjwlr
IIDyuSfHg8W/hBJUvZ9TFP76E3UhOwnq7cSMOuPfFNRdDUF1YHKZwiRbVKEwgNfz
zWJBUZNiVLm9wSCdhIOMcp1NScsFPCcfvjnuKmOzzxCD/c1RZOCxWQueFj5LgMkx
3N1gP0fPZ6d4ANbm5taWppeyYb1OzfHKku0UNgZ8TEBkkaC2IJdivQZe24vXY9NE
UFukcCs8z8sCSocZPXjG/g/UMtIGExvbuCokAoNW/m6w991FhaxWj5M+0FBD2WAT
8QFUvDZ30gdi3qBo3wznjgyVh2Q9FhZCS+Idy5s3teLcXoF2Hr+7Oo4UJj8SS4cy
CIvOy2DHsTSFOAQ4DGeV+9eW0X+rVTG7yLuWxT2CcMrhMmKxHmxAl/RJR7RwYmuV
zB9bNhkURrv/R1p0mvucAv1ZJmiD0vwPRfjKbLjI7PqRTgnVJ+hXkziPnTG9KKIU
i582NPixNCf7baEV4ToY7+h6r/0sc2oBOaoaq+6U8hr8bJZufVbCobvPbaRcojbi
B1I8Gt8ZHywE4pAty8/OGURnmAMcS9Tfw+zROrjM8KUCENNeNhXJN/+wCzsKrb4h
KgoaP8ND7bUu78EBExwCpXahABtVKKZCon2h4Te0hdHBDMSnLEzX47yHRIFnFb4B
iv+Rd+4wtZg0dsTYEvAr9nlx8VfzbgnuJ4RIsw+M4bV1cG6Qrm7sKYxXQsBtVnit
4vEI4Yz9zVQ+y9KFHRT7Bg/i6IH40l638gbsnAE37tLwWKPkiFcfjp/JxSd6FYej
P6vtYpQhxB189atEJWA8807i99zJiNib+UITZkeGBbfsjwmorHCQhr6zL3BF4NYx
rd1LYU0LZzxm3Ulf5yuiaa5djC8xL1VY6X+/aXIp6LchbIjMbBI4mQyVAQeCAQtG
XLrukzkFaOF7Ote85caBRWNivDJt+ws+FX7AVsT/RW6B/cFfAMw2PlmM6PNCBjdH
znv+gYo0ov+wsUtmyuflXRpwTvbtWokbRGT5a8CP8+2cPBe0OhPpmEsrMCBsgKkr
lE97DdXk7aAJQd8ejytjmX0uHn65jAGjvYlzvSzwrCW4LWEIEP/aI2oqYefsZteL
N85s0ZEQyhHgI7IVyPutlvIIRd0LHj8kYLmlkjYg3bRTDJg9jvoAmW6fgG/V0jEk
rng4dUtnYoBXg1+jrEIxMHAJ5KR6T5skxLQQGAwz7AyXzVPKw1PhcYgawGdRaWBd
sYkcNOlKP7unQNCqh1QGtLiBIIJDUQZRNQah1b6WxcRDep0PgSdrS/FTafT7MSxU
yAUrlUCq5RjJlK4rwyhUeg2fNX6zX+od1VltEtACrGg2G6KXmu6mrf/GhFMeSQ+D
9FJvD1XWE065RshyJ4CWMfhJeISD82WqlGIdC0EpR8YuwqTe0o30deDeHuX3XbFj
io/QC6ydX+JekCcvztwqSnHKfBhlloecUDFVr7ArVvd7nexC3q9z3rq91tS/a91g
y0aIekiTNysSIdJv+5SzZMTxLhNi+wLJ0Mhsvu+ZKhAFSSLbw+h8/dfmy/WZAeuH
4W9oen+UvHdimpTWqGXihqAPmr/6i8qUILqA4WUAnFfwMbjtmSurKbIIIXaLoUKs
RjVcTiaUMR7xCf+EKCzAz9TsdvTB7OkJvYxbJt8kW0O6RjzsVQ9V1AZf5W/dmgMv
4Yws+4frJpaT7111Jy9VyfhR1abK/3oyyK35NRSeFAQreqGcBJX0M24/Euwz/wpd
xJX3ChboP+dTn6F/k5MG/M7fo5Mb619zZDxLGs1P6plQuTZfS3S8Jr51GKdbI7uU
TUornopKnFoHytXFoHALy9HUF+PWAX5tJYk1+HI97Q88S4XdYIU4Z6uefbV1VeOi
QwgiuMuuEMxUwuX4G3jUJk8eav5CXBig8Z0GY60qfvtbzoi9jCxkNIhFIf/NqHKe
uGMmFLN4xuLHIArYU909vD3AUFlpxodc6/hYqHKOsVp+BDFdQjH1U6qWsF3L+l9o
tfVTBQo0Dc3iU2bNt68BZfaTKYRsUXhq7aJIBD0O38ieNWPOQlBQQIYRk+xqeHK2
qqArlc6s11QRY+O1PEQR4CR8oA2ms5FVhkK6HXGWWcDUt20pBT3FudE9ReneMyu4
p+LBOVoyLWM/Eh5bME9RuNJBI/ui+QnFvRg9UMgSiQEi5RFxBVWS1Da0JbGQ5kV7
yuSsRQ8FbvK9gcI8KbfO28A9QP1XqwI9+Iv3sFlN81Elfq/PGrRqtXYFgs4ERfvk
hu7MecIHLDX2Bt8HktdgmlUvRvxcOom+/5Wt4P2kwnpHUZRDe2m0nx/VazPLbhaz
UZB46GaA4JVvydy/iC7Xmg+6MUCrx6/uwQyybjfqRQKVctUuAh0/cn/D4l900HAD
p3Bd/ftEJc0OHKfhinKEo1o4rdn/NhY2kpxJ5qC2Ts1PnPemde8aYvNKs/ekLsxn
nzoGFqMO8AuKIgOgJvWbm+8wdMlLW3bQNnXP6YdMdZBBjmVH/tp0Jv/TKJY1syvk
ejMhQWpz+g3/R2WV6SVuW20L9sL5fig6vaa/hmSalC+yOinGozS0FB/A2U36jT+O
RE5ofCURFvjgjnpBA8htezxLli5fOHh1+hZMJxudaa2y9QBt3b7Wvb+2ZhAKr4UQ
UH7fwHgbm2HBz86lFF1ibtmIhyC3aSHXnBXFQ7GbzoR/vAO/J0DEk9arfunPeG4K
YeJW0ExsEcMDrByo0ahpWHjLEqfCCs4RT7gASlDajwaU62MeWQLh348NK35IcoIp
Jol9/Xh1sUPLhQzaw/62rYcSyvFy2M6mHKlWnbrbO+AQXqaUAFJjpN5SRtneEuML
7qgcMvyxeWy7kzOyGp0dvvPT7ofg0bkGJ17k0aXPWQK4ysypormvY67a3tTGJlXJ
AYOvOapwnA3mj+5CsmYtuJnPdRGXZyTWcWL6a0dm+PmBvV8Z9e6BipgKWP9m4SFg
3SF+7U4cu3lrdpM3YaSjRGDjE1TuxG8BxJopMCVlL2lEfPxJTJ0FkL6RJ//U9lfs
JXteFvoKN2321gM03OCPTUborGPVBQ5heMZj/fFp1rEfh0dPZg3p2CGY/mXOpS5e
cxHHOo6wJY6ZhdODp73WmxgDZiMst1+kPSM/xDesYik3Nyf/yq0VrSr+oywDuRL4
EVBhLBkm61oncb3QqIBMgpEw4d65rbZhC8EYKdX0kXHPPHHkuzcDFYtCfHcmhx6H
zyiAcHLW8zStGPqNPxAp3hvD9dEe44g9sdYQ0fTXAPNPIjmMyYAOUVaHGeR1FkQ9
2NmEWgP9MwcxS7QmXBDPw8ltC2rgBRVNdSkRf6xVmxbfU419Zvetq6d0T0t3h27n
Qk8zv+JFFcOxxsixL6XtfQ31xqG9mlpE1Lz/UNIrJFp1XKD6uXdwJozQpPylfla1
zpQEB/Df3whWcSwEfp23mFP8Gm8ea6o7kAoUEaERFLYJA2HKEbNSG6IvTojxone1
06sHMtZWmczPx16k7U3jwr602QwP9MJZq7zdgpymygg9cz6Ln7W15LtKHpGIFp0c
XrZf+hdG+JkkxCkNcSQuJEKMusFk7lEF4lASBctABSvQNxqUbRGLcLju6R4DDmCb
x6dC1Y3HachGa7n9VbyWATUY+RHozWk5biNDcN6iGjGEIlczsmMVvERh0CoJ580Q
bh2PX5UNBkmPj9asikqBBN/TAlHW6DutWxrVUlv/enzXWifndrht4sFwhvsvWxiQ
TylVkmBFwJzl52VJkqXf6RZ024isiAlzO0QYQNknyU4CX+eP5K0XwAqE4pKf2+FM
f486A164Z7kSkrGXbekkeuEsQURRH0TmSHC3kGbLmNP/xCmhG+Vo/y2rAJtVt9CI
8Gtt2fyI8jFqXAgVfk3x2YhC6yYvx5nQ57mI6GgjRChi96pAiTSCcIYkVDgh8jhV
AseuuFEXAxsZ0Nai+MDdvI//hl8eM4G+jd0h0paWSctcCpwwXifgiTNnd11QzfkT
AXowtgIdy5JqGVHbTmfdxdsMYS0ifjPAbtvjMyDdCCFIgKR6snvZyLRkNmfdcTAA
Tp1FLWJpGZ2YuBQ7btSeIisHj1WpsRpH6SsfSYLXj/mctdkFDJfJtyHoUI4FiEFI
B0og02bwm71Q7+xs23o/hLrK0arENxBaZ6OsdJNOhVxe581kDDK5Znf4Y7a6+NOU
hFv60bllfSWCXDYLA6rxmh7QdnWhgMfGvA/9sBlHs2KdMDhi7mCpopBjPJD97bVd
38mUKDtUhT10kWTkbKrOurAX0q2NolmWlwEmFEuoBY5DBj1rc4RTnonT1ZjzeDux
u+dLgXK3BZDYG5hzzFuGygyDW0P20Bjk/c8DULlGgXzUcsotsqEEJKRJIXHjSiCx
G0FpkWCzNmJsTMrp8exh8s/64wWqmiCv2NCZgwypGYCf2Ci7WSgGb+RmFvH0J/bb
PdaV2hZyKAFmxE6gi9AOZgd28cPr4MDD2p0KgH21kOTIN73e+wcjwkhJD9NtNi7G
quAhAqTM4rd+7svvt/Ly6iqaTsbbzWPEdRDlIjsquklJHd1c5UdKYvafy7iecYYq
zIDknkqy+1hp8QHuEC8k/fI19M/uQZj0MYS85yWOVtoYFf5ptBfU9ugD7+D2NI9U
juZcmnBNwdYThCBZNWKAHrYkXbCbYdXaPwFZV1E/udDYLlrhdyVa+DahGImATLm1
OzNT3bNWSId3gz6/E/+vlEhRU5NyEGMYRW+d9ga2XrprEhsVxErE8fXzp/jfegfK
YNgp765e87R+HOxaJVOtRfS1WyQlfvdqJRlyCVgX5AvWZTyL6lVX8mw6h2vAGiTm
Uftw6q6MJU7VppyrPEYwcNnT+Mg4hMXuFve6zLW3jqSWMSVm7EYIDOT2o1JPx+1p
koEVKd7JgS3ik6lwgvm3kEmYOtExCmokx0Nxsci9UZ8Xe/6KSK0GkuoUKfKfxntL
i4tCgapLDI/VXbnhWIJ109tvkqM8NEFn/BGPnPkO48mQrSXLrqv4YwDuMA9iTJd5
85lfcV3YEfLOrZXfMcFXc+T9SdBk4BMiML0XXnHj453dmZnOnjyu04RSBLIx1svM
pzZNSUuOk6WZtOWQoGxBqk+vZaNaFESjg76qsJCy1k0nmWSwcNUUnZcSneBq73ur
s5C13pWKxVBwpzP30WEYzbDm2gzetOKt5Y2uv39Qsc5VO746sH2ThlIhqgVgfRSy
RkBw4IJboK0GpZzdG/nJmm+TP228nXF9g0Mktz3x3LOCJll8Ltmo3Qn48/CuUzNN
okVPO2EEyNMD3HPovvl1fw1SY/vT8pFRWcSSO8QLoYHhpcL0orevN8/mjFAHyunp
ZDBqXXxrNBfSl4nEZFtfp5e32JUyb3Lty0Ivju1c76oa8G6M7DnG3YPAk3TDiQ67
1Y3qwZtgHuKUkncdJl8TxQklt6PaM97GEabv6efAGfDFOQQQDbUDddsms+fI4pmu
2B7nAU921FU0zqohI7r4gxmBP7i31mZfPDdcFdfy7evRB+1Lx3GCOR9QekAQsNWq
3zXmOcO0G/wKXBvQa0DPFwDx0ObugAs3gHElEosaetS+RMF79Ygkc+2OofjNOdAa
Fkn18dxV8MxNJlxBBd4FvqrxGz4tHbE5yS0hAQDV60tk49h8kvjs/uwG6mcE90qD
5HvsJdGtTj6Iz4eyd5nBdNV/6mGqpumXnWSB1dIkxS/iIAArDfNlMIiqFAynqHom
TdKfVdid+b2n437PHv2SdwNsB7OfECoprUWCNgfXJI0Kftr8uYpBGSkJkWg9ftSW
4P/IV80iWRC09jYqyiFaPSpcGGEpBKkZM4UBW9IUUKy9LUZw5U9BbX6Qp4Ltd1IR
rs50JAuj4KdmIkhQ/QvwTDzN3N7EXsQRXTVhAa0pMU9hJVcLnpD7n08BRf7ZtZp1
RhioRRreNBRr4JXhxKuTkqCpOXxg1VHj9MmEpr7+fRTT2CdOjnZpZOXg67nFjFeW
b6acFpUIv0Jqmz+gV/KiOSed6aF4JNkyiXFyHJSU7homP5V1K2+D0472Q3UrJs7f
n+Ru//kqhibQGv7XPOHTW9RitNumAaudlrKLnuQqadI/cAuMq/W0bU3+UAfqNL61
9X+66K3tbQzXZfBCDmPrkLobCx3+v2v4MwiZu/CujVwyZ6Rht91aKFH/gdV0qSF2
KlaiDgaS6SLypl1YKMmI5C5MiyG4zIrMHU6h7f3oQ9PjVvWyxaww0oY5yFdz6fVV
gFLNxMw7xYg4woPhA/kTxCRoclAhY4jN+a0RKn/8zKWm6oeT3opIzFT/n7fdirT9
UrTkxg9+cOJ9kaMAK6k1fhKd3jUtJOZ6BLwC+LN4959nscJ78yEsYCWvFG/vN91X
11CRqjkw6OapXWSXG5Xw2WYK1uRHj4f/6Y/znxk/MXXy2LxbFWbayrKKH1hIBgfC
7uu4IX+8O1xhb1pnuOrCWIT50EidqEqoolqPAxbe5hQjNPHASIsbMspEHI6EN1gH
H2lHzeXlm/CkidIhaYeII8PrDYvLPmkOUBkl3QnXIqK57xghrmre+8KrH5Dyf7kC
85Zx5t4NoT/taPNdUNHig2eeLbtgIIIuYrvHG5nGi4CO8GcFKzcGrzDfK9KpgDPs
e6+FyF366pAsy0iTYUrDemb3/NMV7Qj9jKm/RPxpxHo6egyO2C5HYHATOZFRG/gl
UPzXunYUdfZeQZ22w/yMoVVP3mux731GfpgWvDXpUlSjKz0WJNHolHoJ/5dphn5n
J/k/E1yLQa4VqjMH07HEXJ5GCzge49va+UCIbrQXy1WEbU3EuoDggWKg7xpDRmxl
jWdjP+esR8+wk/DpiNOX5ieGFpU9BRIM3MeldoPBKoZLrHk72Y8UG8gAmRMs97r2
GaOwF05D/ysnsVUXhnUneGNqhEq8fomSTclpAzQUcz6lm98boCFFki8WvHOjHHPb
EP6yYlaFh2jFI6cdvwyBWGPqrJ0KM2cBLdmpxT9QzFb0rzBi0mXe8DHxQtHBBUSL
Vj/iYR8ObvhOWLWRjXPV31bCw9zvbTb4HMgnZWXOcT/a/445k58Qfj28N3NsPmnd
lhfQh7hIjH1i1BE+ZRgIrMyl0kr9UfMAMGy4SWbs9iT3wCNyPumVa1uWEZ6oXUXq
gkyjl1gGpq0l7wJn7HQ3iufgi7aaXYi1EdG+S0R6Q05aB8c7ozJ6pEbTZ9SxbzY0
xynGTpRFClGJ4XSfM6HheBiBiZSU1MCoEl9KRRCwRowYY48z97hW4w3aWENGbkM+
+mPV0sVXyHih/XCV6BNfkQWzkSBGH4fAop7iZgusWlUpHwyzqZjfOPH454IJguNB
3JZJmkiyljAkKIwXNYsFRUQ/KZmF+do9SRtgM8QLntmVXdTdAJvAJql41R7TH/py
bmcYmF8HVn/FRmfrniBwY2mDdMAXi4Fzc/ZLD71gRSRx3mDNMiQUnep1VkcUpmpd
l5MNj6LbUcc/BNfMgyPglMckPtn5ktS3xdQ6sNeas/BXEcms0BCc4TNSYRVwXKUN
w2MFouAng7uVMqIdwOctIMJg9Z+xZIsJ2TwTzDRrpbXNjDARU8rIxQYXhpdnP0Ob
EiXmG9ffbQ4pMYAJpMqfKcvjQcZlyheN3In1EwPuayzIiXm3nt7Xt/nxvokMPGId
fGomOu5P7GVFjstn8iSio9GTwoiXpMf6sd0YYv2WnU+M8NXiXxAs8sOQlEKxDKmL
iAW1EiH/ba5wB/QrNrQmwYdqBT6Q7LoaOx9ocfjU7a12XZ5A5pnQLnPgTQf8UUdR
t/hTlxJMEPktlYouqkkaR1ZJjvIznrgZQERwIi0g0fKU1JzU3HwQ9XKlBO+PDkX5
cyUdOyLXAlcKICtcDio4reIg6ewxxxt/gxFpWbVl5t/6FExsnWkGos9DczF6LxFz
wHBuSjBjpTSFMnpVRDpHRczHXUXdQl85ch7IAOEjebM91+CmOucUJTl65gSssVgL
VKVwN+HQVv6oqgapi5m2H+YqRyKqjCNy/TMDIQE30R6R/t/1xA/WWmKf2+ZLajUl
l7ZXrWZrJ62Z/OmxikuHCUchJX5Lz8FERf9dW4Acw1cxQzY8+ASvUeK1rL9VT5YD
GvI1N2W32J9l6QRG+V3ykMA3rE2k4z+E7FZuFE/40lkk98bP2T9troofsXb0hGsq
9qCHJXlXR1hfvE/rd6gEulqBh5Gd/t/woE+dhOccc4PS7niWwlXr9SH71B/f7n24
vVlUBs/lltZOOeso6ScPbuekGu8snpDtOi0vkrGE5Md9V/6+fhSpUXOGtBwC1JzW
e+4NVJ0okH0ZdhcfJyCTxswvcXbYpzYUWksLR4IX9cZX76weOaBVpg0ibejGbM6E
TxxUEl6Yzb1fd3EU/5+bidIr1MfEJZrKPRNBft9pFO0h9odd0Cg0ijownd9OC6EF
UNM1lBUSVM5AFthWy0isGs7s1N084fkopBDbe6cAlh60VX/HNLUHzcaU+xYTWWZa
gLH7WFSncQ9H6MGrqPAcf3SwcVZeJZ9+cqvG4v0iotftZu82DfuCEBpBsugwfaEo
gtv1/lj7NnxE7b/KrQQcj/fGB1SVM+r6XHN0Msuwd5NgsNzgvQJTgAmlSWajDito
sdXJw3MGnvTCG3mI58pZDqtKchDnYDvFHYSPYvohx4qNIrPXGG/cAwFyYhvcCko5
X4sqBLPmnPvQ8nWSJcug5uUQq4gFgEQnpuSV++ZzalAAkdB3j7cDlQR8CSL/HKSC
WWf2dyBRmeCL1S5D0+SkWc5wdQpUSQ19Ms+4aSpWQ8sgKiPxLkI6zah6gww9ATEi
rDjgJ6fNku8yihLUZBBDtleZS5OsPzDUD6Fi9wpCQIzKcOh/rAW6VvZs9IuqXzco
3FUyEfqI2ghXGChivYv0Xavckis/ge380mxq90RSK1F+UAo/kkhnXZXanbh2C/D5
xc+DwByVaQl2Gz8LX/sWTBzHgT/r2orA3wJPMOM8R1Kvr1eAyBl+zR/ahzht34Ev
7dXNTck9+81OQEYO9KjLsUJGizVPy7NHkO+8+DDW4pbbZs34Ok2FpkNd5IQiTSgZ
flvx24E3YyzRJFPs1mChQZ/RcJN2j1gxCZSkMbKoNsBq1E+M4l0ovQnEk1DrGytK
y/iBkjf1/bvv7DbSkUTHf/HQSxo3lrRag7wU2R/3c1CTfJKnUMlTr8ujNS/3TO5A
OsDbUfh0O302d+fQSSal7mMKFpber+y8N3yoqkudJsWRR5QAI1NHAlD+8hYGflw9
CHV4yIbtUE1JTNCU5oN/emhfIRH3rjCMtHoCGrjpPLry0TVb5beb1NzX7wpOPcMq
VKcrF75pYOSH+TP5Cs+CV1G3YZUplGfefHksQY3ohoW+0tgo+iYKFn+4IoW8Kdt5
nKYETvu9byM6pqfGskrHi4HjtVKxNCdzXJlJwszSjW+xBUCXE3clZC/fUvdbqo93
L609oXq6FbxD2rD4BAQWlUe/cSocFiZsYo5gNz7o0poiHZST8hivIr4t9zEqgSnU
MuTHQHfCvIHuTypgT4Byfzkduh8Ygzj7RThmoMmUx56TGJv1IQ7tOKQvEDcLVo1h
ubLxHnHeeYREuQ8D2Su2b8TbBd8dt3j5+aO5719Qofk3trZ5M1nDV5CCD1rEXrSW
dpXom3YYjscfNLjce/bLioX6HW3OuBFpDPhDAh9VqUJ1+Wa4dBD76juqH9zr4Ltp
L+KiplVd4++S5MZW6KXSwr6vDrPHsJmc5lcazBvkFNZVExe3WOGB3viLXTGhj4vF
H79siOsaU3e2wITuvuIBgss2YaMV7RE/ZkN65HUVqtUFS/tCfxFQMlncZNJl9ZxM
zDW/HirISgpgDeYuzU3MjTiN4QqM+yghfY5HFAYtOiZTGPjrzATBXaMX0CDwcoxe
uB6HFIr6EBrUy8KD8hFx2UEy2Wg97jVRTMumegPU9QO/OhfDslY5aH4/SAL5zM3J
P8QFxcyZNRXF3mn8cDkUwizKw8ZmjXfHr9zcoDgQAdKiNtvVpX4TkGTChwzUQ+5W
qI4dnvGLpTOJ05l9jws83yuYrtN9Nc36Am973mGaZsZtSBjxA5HTCQHfSCzxbSZZ
wuSvaI0r6aq1u7R2dVbACD89NI0i3FcYjb67QJ8D9HKZ7F7jo4cKCSYABXupmP0Y
XMv0Vr8ZQO1iv5oV5sUngViSP0qzYTLMDMZjflIFYr2kvUVPALzUz88sBqmcmyqY
zWmo1lauX3ejvkOrV6ufBo4pOmJ8Zrgqkp6QrJgCjvUoFt2ssUn/gNihs2H0pTdv
dqVUNDhc3aSqnLxU4l6KOieu/lUww0n9qf3txD9hSXrBpqXt6K4RG9t0XPYgrXBC
JoHzMA7EKFcVJtKpKvllark7zol499A6oUXFbsGORiU+3LciEOGhFCIj3rnSdjVk
N2PU8oWzV25LITGUNOke27bTZGgbFqRHeIDzOQq50tqqH0IvPcenEqBi46e3grqo
vEPt7Lb9Ar8tdl87/GRW7VTVJiKJ95VOXvGikOm5KhsyRV0gIzLC5LKxtj/hHZOx
eMpkncbsrz7BEIc+nQqulz3qr4oK3cM0yxzKWiXn37Uzwuvx6oM4KCHejHFhW66W
Cgcxwsu3QuLuqftizKZgjkgmvKbu/OmjrzW8Us9DIm24nqNYYy7aBzZZ+0NpRZ2O
F0StNExktHicyqAdG+tCO71SGDUY67iH7NVJ+4+3pqeLx7wy4dCQLk+96Omdsb/y
0PwuPoDoZAwx1T2J8L1uKnNISveZt3ODXG8XduVx3rOx5YS3LHtZUPoAYBKZ969i
4ODneYYelzQZwr+Jq3Zx3oU59vmD+Tamg+Mxu2C5mzvoIV6LLN+zEvRfBAeV913E
/G+eaHhiEMtab5j+SctPTPtF/+JCh0pEYbXvkaH3m8WJTlvOiUQ89pe9EsSEoSJy
7WkQZZDjFX6M51cuOd7NX09I5Allh9vh+c1RKrN8XfzONQoJmhY2TU8iiMCpatGE
zq0TrAYradkVqs5KpYyJFj/kbd7lfP7Ya1cc+S4qvaq2qR2p39O0TRE8qr6d1THo
0H0vrM9DyiWeIlwZkHCbJtRuv4TrEv8dxEWoPlkQgY8T8MRehpaHD6GIAYg2Z6a7
aR/iM/lDeBtM4+XtmZvsRhhQbP0ETgk+2ModOH5A2/Im1vM3WwguoM3bqJtvQQN+
X/TlgDbRXgfv+m0Mmqdf13S/mAKcWjzrZGjfv36g1wnuNv80nTp/UWsWyiqcX7k7
YfCJYLlzTkykaS2aMmRC3Sd3ILFHF1P/gFRFoAFEhfQX2ZKIY3wB6TSxk142UHdI
jy0rpqptaB/sKlXcr7hTwk36scXY9f+c0tKTKz9uX9/wf2MsYRI3SCddrbjUBHw4
xLcJMuPnMbZECRpDRa4H7uUJ4Ivv8jKh3IdOwZoenwhNThmnMjm1EWl4MAWDzfqQ
N98CmAi8GVHfNa9Ru1dAkxueIjlR2NjhJyBm4AYsxNzBB2PXXFtjmY/AfO7CG7id
sltWBWMqi6Hf85SOSiJtJFOVfBt+cYqEfg5PTiMWbm1srXCfgoxhuQGAhWguZeXG
H7CpZj9FnFasnTw3eML9xsVNajNAXG7VzHlciOLvp/Nl9rP98IiZiFm4Ijo8pWWR
oIJOGZEp19KpMrSqt04w2RfJY3Pj1TK5OCwVnwxYVpldCXpFjmBe17+nzT7Tkw/M
jtlyUBII5QJJUY4xpwEKcRZC1a4msrhSS7eB+HMNUDH1Zes7JJe+r/ZkvkAHL22S
g4+8Vn8CLe5BMmBqiF+nmLDYYSuBXaiPpLuRp4keof0uQ/2EkuvF/EHA2y0m/SZH
UmzTIVurmKm9Lk2wNz0YffUan9Qsxn2Ed9ryMVyLm82utpHge6XFjpqnIUKKQVtY
nrPWgmZju98wEn9Y528Q3oTJQT+dcFWUXtRY9+Q7ylCwg9QhjRisnDpGQZViadt/
rNnXfAK2bptQcOKGa6V4uQd1J/mUlUwHidI7NtzoHDan3OChsJ2CsWZdPEw/gRQN
gxDV1+pyLOCZ9Vt39ZQbPc676iYx9AHUvvY4VWR60fV0Bmo9QXVF4RqFVzlO/fXs
0xFdLU3p0JwwD2uXA25A3GsoWvWnUpdCUt2s226KvKAb7mf3r7bj/vazG4Oz0ixg
rd5MzS+YPTBWhYi8NlNJiYM1fUEhMlNf3OWxkUgt2I31+wJfF70MuES/pciBjzI5
z53qaL2cjt0hehMZPWAOAsEL5Mg/KbdRFMX4WYO/1QczG1uLLNQMIolPbdpvQEbY
6xIFQvoxnB5GnTcxTEum8GlC1l/8OduOUgW655+appFZfxO9cioCTz+bCqqbcCmi
vCsjOKg9cb7zY3l+yX73yAzYQWnva8JH7P0yCjKFB2WmryfbPsLtblihwfUYXr65
GCOpS/I3WTKP/BbYHr99EdotIr/UD5Ehl8OnBxcb1NZO8pZXl/xZxfdqKiMSd0HU
ftgVTrae+ZvdkCrDkqiOjU/QaqdgljKJmUGV6y4p4+DlQAlxPaxhT/ZwWsjH7kXl
hXuuqEjNGyv8aFs0gKrC15Yl8s5Uo25uJrW14FvLERqCyqGvu6vFnaIy55HJmccI
40jhlC8owJa1wcNO0yKpLLeIEiqYRYu4Bb0wLn+FNHcQ/8Pbj89his2PEl+i1xkX
HlmegnPi5Duls8uMxFN1sldyuTGVnZLIY1+X9wxm11MVnHp6MdTOu/Alrn6cuWxq
LwbQkwBjqHULcweyeectyX7FNUa7QZwtL9vdTNGpz54fPgPi/VmVZXAq+6L9eV3B
JbHOIGJLiasaT9rpZXu7T5HnDRuCy7PXtJbn8vkecAfN0jXYLM97Jd+6bzymjAUG
4OYNb/10TxnVH/TjSXt/y4H8i7u6lh4oNdQn8ivvV5DIY/jXWBUEecWh7B4WP77P
aO2WPTWlSf29eZ6ksYHt2OjzIXmLCDWwDHULX5ZgvVMeCTT18ZPPYcs+LTMXdrQF
fZPgKkGFXp6x2aajThT+Q8qQT651bbhe8lDiqt6/avbY5FivlWSM0Xj1RBNNBGsu
c9K06M5ztlQvlhAhzyfDHIH6m5EsJ/KvugE84jQ8S3XDr2PtVbilNpItbLHJMa9U
r6RalvtLrvqcgCRATf+khYMkDvAtwUY+iH773985iQKULJJ8rhpCwUzhyzvmcXye
Ygm0C8StZqV1PlWNllQeCMs9BsnEFJYTV6PgbiFn0R95tf7jao3La1rLEMXE2bQ6
XzJnlvABxLYEKnsJUh3Icz0QcpgkdVyGijzxJapwDrxIz52TUyhLrk/kE5AXyQnu
rCxwpLvw3eHck5Pnbq2QUhrKCOsvguiUNV+b5cI5Qah1eSob0WL0iH9FQE7W7MDz
7OOViIB0wle4XegyWk60b/4Xog/xAqtsBQYcyKJe29LDWrD/pUQtmxsjFsgVrl+v
mNv2TBpOQyXm2bafqv7NOEc5t0sCn74l+ijXMRO0Q9fboJC6djO1FMjHHv0YPss3
PVb7WdSngL1BaS85/T8xstJPnAqFoDQ7+Ls9DSQisb1C8Dz2Xq30b3Ped9ysdO9A
ma7HN1A8O9PHWhqJ7TCNzYQ1HgiLI5Iag/4QE0NL1ihkt/K2gh7vbZWcEwCpe4up
CKI1Sa3I2VL0MnnkH2vsOKNWtRpi126AMrkm485t1HHSohgVvH4UgnyR2zGdIJPQ
DXEQbgIMOZMeyokTkvo8HGdx1ruSEukE1lQFN5j19NGu/3OHhx8GE+pukJoZCVzs
ppLdI/n1iTkyaciT1aw8oA8o1IXSepHGuhq6S7dZdrjS0S3J4dpmlL512fSwPVuf
/op6eJvSveGeSVdAnkKZp9vBm0R2inMznuk81Q+PeGO65/U3+OQBa/z9MHEgFwKA
gG1cBnD6ypyVa4ymhNLvFvZfTjUshfWqi9i8ZvQFWD7ete3Pl4s1Wb7EmGZiYKcX
f9h87piXAVn8294Xq09QhgytX3syLutcQS53eFekX2a0D4spdj2rGWUE8j1FIv4K
VB+HPSEUy2yxjxKh2beViL4ZCe5lJ6yeYZWP49nQoaBUl0+vLXXJxqreiRGpnZwt
WDS4Gq6ZqFeJXOz69ayOI3h8DLFrzdEJy5b8NJdVpYZGOBwIWjcfXANYp+yRjxT2
KWAXR8RQSeLTfRNA+9vimba0i+eASJBxeixLFuCTmIbGQiPHuRYmaegIxvX4yQ1L
5gzjffF8lthZ50oA1DdeiGOBBrsBvWj3AI/UwFO7V4lpW8XM52bDAOaR/H3zKhc5
Oz2TuzFTNpckkSXtYyveziS15bbof+6JRUrby+sIQmunelzh+j8kj9EOuKIPl7YO
ygDJGuAyKZYTDSlyBU56XvL+GVcF73u3C5P6SdRceO/YOo/0stA+80qNprYrTFIW
0jMYJsbaRjteXmv47h7IyF3U7Jag54Q119diyAOPAs/V68JMZ9N4TGJQZEP2yYXY
UUNhkDmz20X8yJjZg6P/sLS39+QWtrXMmxX+Y6LQWJBby8CuxA5ThiIlIySRO8q/
J01WM35Qh7D5VFZ0E3AzXmC2DOHegoRcET/UHv/qofLiwSu2jQK/dDzHQ13XmZ71
gvwyPpYVGRsGux3dl8KwP7uCOwFKqXULGam8phzEra0T/1BUwt67mMCNo8IeZRJv
NjNLtACZy03opSPQRIeYirQXsQR/hebQU62GeVMTgSU0FNCZGgZ3d1v5rhvFDcSn
XxJ7USHpR5Alk2TazZGNIq7I9cPSr8dIPnglS8CqRkYSgpXT08XMX+cwzxtm6/JC
hiSPhMlQTXJPYDJqiRD3V539YbS7g1bDFbig/6bvmx0Bt23ttxka2jjqNotg8s/9
qi5kLUVCHglen3pOS8StgG7FrgYbJ2HtY90hMBkodHYbMFpMsSpwa0mSJD4aNj3V
PiLOP2r2nrt4mwlwZaLr6oLRbXIULMrwGTr81TV5ehTYxjcKbYSSLMnvea+T0TGj
3Kj79ds6nkQV6RznKQ5uXAXn8FSNE02lhg3sxmqyFZ7P/X1UegH28SdZN1zLlYbT
o0f9MJ6qs5NmDLMcmkEHpPPB0PK5IkLR8oYJM8XgUUHykAHk8xJz0GjEUvO3qapo
2n0sU3dfNsFavKocJC8CA43r6pOtUTwQBm33kn/kJPk7bfyhu9REzE53GdGDvhVT
hw2JkQeiSzzkqrmvrIhjPXbfETZSC+LpIFWaWgfWMs1AtXKzvEAsm5FEE/Ys5Btg
Cd6psqAgO3abOGTKicNtfWEXw0U22XeQZO2jBdlEz6xnFYVQNQCTGXaY+Xa7lv4M
acuKU8pGPiHRHp7U73FY+GQ28OxjywTsbkaFqDu6zS5nXVNSlXXNJOLBMM61GuuX
/YRy5ge/fLGhQTGCxxM5tfnvzYxYjDs3TYKr5JL+3QrWjBn/Gg+pnsAZi05X2Rax
TJOVQ+vqRnSCxKYh7W3WL5cstemCj23C/Vt9unj8H8C8wcTvi1c98lF99QGelGpv
tNH6TVmtFzJ6yEkXfK3I5J8QGtcu7rLpFwdnKdCdlWU3HuMewclsK+dYzDRXd/32
F3Nb9MJ3/kJkPOIkBtZu0sEoAqJ5Q9zGrfBlVWxFEQd1zf21ZvIlAosLzzo2+1T+
GHv0f4dDQii7gRagExRPEsnwGopt9SkU/nHGlNpKcV62u/EplXaqtgdbdytV/Tx0
xJyavpHJI4x/G0NwqA1q3CTktyodTOit/qTTZuMDun3UfuqSQQ9sv6+/AVmIXN1y
boFNOJELLHnjoGNQJVLi6kpcjjFakDTWq8Sy7JT4FXdzpmcZYpCQWL6ynhN9XD/I
v5VkfaWa455ezl5ohfLR5rzSKrcGa/x7Mth7DHijAPcodKbOS4mIgT0n8x36Hhvc
JINWpa8o1MCH7kPO7S6HvlkPNyM8jz5Q2ew3/E1SSRrv5Au+C/Sbpn25ohLTC8Vy
B3PL8Mx3H5q+CSpUV/vr6NQ1owg+JhSPpVcmBa/M2+3VSKaHZP4sF0UBdGqxi0aV
EIUb7kul92KrXNIt7CCpE9OPHcDf0tNxLP7LKeXf/n9jtvOwm6mjnQAgoO2sjR1X
cQczuxsx3IEaD6LAF+BjRFgqtt0Jq3HumOCnVLNUpBLekBXSU0XOQlXaddCCK4LU
qeqkdAi+Qw2YR4qXhtr/IVWU32xH5PphHlc+d5uMMiQ/fLqpgXDtfPiIdepSd/TE
9jfrkXl21XGUPfErpFNVxxclOEdG2rWUJZ6U+qCf1MC+nm9khG06yxpPxJxSJE8Y
kfFs88way4ET9c+ATT/F4nIyPWvf3CcexXI+vTWShV8m0wzF36+fgga/5JwHHvBF
jjodDHG1BsiY3fGXSZNbShDrqWtym/X8J+uO2r8KBjVU5EGS2YczGAHtqYamB/Uj
Az0nezU/JBImqlZAso2ARb7POQYL0nJfBRvAE1VvUBMu0s+ZM+uC6J6vQPwdcZaS
Uw31SHv4ShvPZjXQXtDFm2sbW40oRGYBYPNndta9OJ3xyMVYSSkoHgHmwMyiwTBj
PkrRpnjGHG+yrQQhrjetfMEcXCNzRzX2jFYv7TkSTZ5aLrwVJvIjtGN/p0O59sVt
P5CBkpWiwdgcOMrkL0xTGwNDb7/ANj08Yho/DGts+LS3rRiU2jEHM9cin5TGzBln
xCNZAevq7VcFQhom1jb/5PE+4Km776eBozIqx6C/OF9fzXOEgCr6gp0eMSRi/d3j
QTWiutmmnZy1XbJlc+cgaVx/trXqNsVKoqoqGDs4sYCoAB9cON9LP/A1J7L2u7dX
YyQkfIr+JtxbP2AXXbYsHC+8Kn2OIuwSQvIItEhcuYqUnvm/yNF+VupNh5YwAbX4
V0ALlZc1TYEQwQ2+4UERCNuUyw5xdbMiPvrdWDGMsQFKzhRRrxcEGRBZlPrrwdBl
bJybScePSarc8HhG1JnLh74l8nuIkNPLimOGqjEfdqrORhS+IrjuTtH90boZnpWa
XazGW30Pkot4WWSLD8aOno/v/OyotjZdClwPzRm+1xEPxtQMKdhQDmab8naET2zq
1lf2ozkGt1h/tC+4WpOYaXJ0oUm4HzxeM4GHKeVHGJmwFODhS6RAU/AJkci4Lpnb
2vlkH7yNB5Ny+XU0FQFemsk132Vbolrutm0dJRjrrVpdpEKpWGP7j2IVn17qiT82
8AnnmPaL98hEur6vntx5yjCU9ZT+RrrH9sTfPf0Dkmz9pWkm7vSwmjQ+GrSKs4Gm
rg7Pk1/Q3cIV1Lmkm0O3icXkFbEXTrm3529BU369iE/B1n4e472wWezXmypkFxDh
G6NWhQ64YXdkrWaAkb6i3QJ6a5yoPX6XSyTzdZLbRHuuEvlDuYcNQs3sCyISxNtY
8Vr3w7MuP/IMpGWOYqi1YigPsr1nLrCaM2zIo4d8sxifF6jgQvFU9LVXe3H5DWPS
WYBOolFb1exbqa8lVVYdifAzE6+c8/BoRoI2Me7uwdKDi/pvfJsekrpvsaRFzwlv
VdDUgnQ5nQPsxN22HNfA7F/aGeIxnQkBTjq4LuPVavpcZD9PZN8HciF6QQ8H1Vqd
UdMPkEZyNzsBRFPSb7CRaMmmU4fjBu2DIMmV8Ntb6FElQ83vd82Y+0uxf4grfBmS
rb7ybscHjiw6/woY0nF+q/vTs8U1zAgm930us7bq8vSemc+2cRZknkRgPqrFrFyY
AFRDa/xvHkR/A2t5XUMmd3S1PCY7EZHdTFencfv75GWyf0GzngI41Z/CogbA1q/M
dw+JNrEYn/oeEhNS/YkaffDZWPLg2h5gg9V2Br3TXGrDhBqZxQnC9vd4iw66iXWH
9zFTmxBwwVVApGsX70DJ5wosY2pFhHu+CnvHIzb37mrzh3gD6GGGZP0kQD3MKzOv
m9gguyLePWpfjRhWhXK0D2Z1G9n8D0j15Zf4Gnmn42ZstDpitGqiPRc49M9V9iNk
ZNrb/DrG13mZEnBqXuVA0Ld4VaeiI0lakYN3Nb5XX0g0QZnPlWoIphfIkXr29969
v5xcuBiqjIRR6HKeJJUY4Rbrd/7mw8d5FNQaXSFNUkUgcyDIN7CQ677Q4scJRJ2q
1GRr66yqZbkxof6D0sY6gypMqNvIK76W9ibC7D9GgbPjgLaRDcgpT5Xp2piyHu49
T69Pj2Y2B4DCACqSEEabXRVz0oew861s17R+k7cMyOQw3hqpEf1zJXW5aeO2RQ3J
olVaOEQrhomKvpwog8LAhZ4LYxqYnylhm+MGTe+Xix8m1x8xqKjzQ6FTRoTuDxbk
XNbZRJc/5BPbniW5N6/M7azHpY0c/V/+UIHK5uqhB8AIU+NJ+oepXCG8K8Bo2FLC
pU5ZRMoZTGt1k+W55rSl31HlDsNtf/LBKRkgyev0L0apIMaWchHjfsoZx0KgYRtO
w7PbJaVgf7ZN15lN7jdCuCgN7TwuFeEhkGUTa0uTzlyraakzw8BcW4DnXlrtpSbM
wPxyhAhbTziwDQG3ra8m54gExMr6CxAmgcvsUbhb/ctxUhY+dCNhgPCuhbrvflG8
kPIl8Fxk+TdA7JXdXf13GpcMrcTmjHujhIGHZZ3eHGsfYmjsRNKomGyWR2BbXizH
AbhhXlAY64XW+XFda2pQR+jAf0EPqbMo3Gbsa7LS8NVKjxreqYrwNmFCedkkwHMN
7NBpPQY/OA2mK/sIne7tyN7v90lRLlSTN16qmK+rdMJU2tNfF2KC3BL9hb9NgCnM
o15due+nG1OhLJ4sUP9pu2WlzfGd4woKCNWZaH4xAjRIRxu8fNYeU2X0mWlmQpY+
9d4d4rtHY+QPEhF9goHGtkR2nXwNYweOGdXre7uWS5BV3TIL88Nc0RTsayKpiuRU
pbCq/iIh1L53gr763S24IKyK5n2pAr7lKOdGZoDIrXFCPAxLJZ1YZZ7SzTlhw646
FuyijaWDd5SD1d/mHbREPr4/2Ob3mKDu6/V4avQgDUuQQvjc9xOHlTNsw4svCyIs
5iFgorvPPOdLBmHru+duu+JNGcDyicgeP12warYtpCBP5mDeWxoEJXhb5SJnSDK8
e6A80v4dMtQ3rvXjTtxbVTqSKV5YYTUAbtOvrufiUiKv6f4h47yKTFSownt24OD2
8gncOl8rYfmyv/FfSvBmS+bfT7RdUpgBv5YpjTYJMY/M4IgQTv2or5lDwMT09I0Z
IOMsiRmZSK+mfM3Xrm+Ek2TMa9bL9L5SjVSQA6cTsOeh+BEJPJqZ1X8J8EJMPDys
T8sZCTcK4wareasRS0a26vkDuMVem/vT1Sb3eZAl1/dafh7ZOd0kD1Rk8hpNPRZR
ZLTx2K1bkeW314QfXQFDLpnenSaPPeFqWhrMboeleOJFS/1fCEHIWLD/2X0hPXAO
uLh9d/1Fw6JYysU7fzhUQb4YtGH6bXQrGJBRB7kvYbZtnCMY44B2IwOAzfNN0riz
/e/5f0C5wJGVj5D4VYZwpx4ZKKx5rNDI6StAXcNBie+3Zj9aZyB6KF4tFkGd3GQz
VSxstdWe31eV026GHyr3Qc2rA8azXoajGWdWyPqpXTYyeWEAS987Qc5iuuB2KaPp
OquBHC7K+m2xPq453TXKm8acllcOvchWjhHiEjqAbAeeZYtnn//FfH6VgGpzr1zB
9Q6OYDq232WsrPG91Mso0cpYnAE8WNZqIYbIpdblyrXBjaj/xZZs/hbokmgi7tbu
No2lhaHe29BZJJcNsGUWPk+0DfuPS0Z5+A8TWJT0CuRO7qTABKWA/X61za4RPy3x
n8ccx50mM9LSysQSAmjNd9bdyTDo3/CY9t9PijZEA3kOTMh6WzUQZN6aVYZZZeIa
GeUUTMLPIcU6vgyuAMwrNrc+ATXXNmyujpeVp/uAYoSX1foQD6fxre0pV3fh8ERy
amk3jJikW8mtXyj066JN/ylUSkRU6TRfq5hpWZVIvzi/WUAbSbP+L2rRmI0V4bZo
nthZXqd1QmNszH/cgpCeam9l6Q3gUQEE7lQ0ZS3OgZwa8e/SErP3dvEPPZcHJ7+w
27Nq9+P00Bk7G+L/KOGvYGKoPqDmyZlsnSxjwQ83z3qZn4TFLf0MqfuLtTqLVb6T
18N1iYGCGM1QHoWU/tgFaaasIoY3EVRTHuWy9dBRncNrlzEmqQabX+TdtNwCCAxU
XuWlt+tV1nqQnf7GGx3o58iOdKYqlrM1c4LvHIYYSslSuOZry3QUrK/UvMYgGPpZ
ExyJ4RvUuW0QdRAr66M3ftUY56YipJdULorrg6nNjmyIlCGWcrdpjNgyOMnIfjoA
z1z/RMLCrwb78HmnOAuKYLdMB8xPVU2nBIhTX1k3iIkCujWDtFGkQkvl75oAc7tB
TMBdCXgDgY699x+mBoyMp6EgRlSH+Xbrn9Iz2MICVQIvZ+E8W1neaGU0Yin1MSLX
sbQMzgUhHLQmHwq7K9/+qKFocah9jJrNynsGqf0jPwAyvcsE6sIreMSEN78aSUuN
FnYVgy/wm5XWYpCZ3BfKWDA6pHxBy076KYcsfhl2cTJe9PAi33VOQ7XGZyKqdcKJ
aCN3fGb0eE+wOrWDFZhfpgdSUM9ePQmh+QhCipdaFqo17Efre6E0puG4jnPSYQ+0
qijHkux7MAKdl/xAxr92XXVf+yLlz1m2tJ99pbrRPQzcMtNcK5bIe0pLcZkxfJ4I
8VJOctH2B4cN/xyVvmXXD1QDX5PqFCbpOlyUD65M5oylGATpU87SOhb+NYaS32/N
SwQQ4yJ4UYte0dj1M8K/B5zFQ91Hx8cGAQECUllqmTOhRB2UuGJhwtCCfInhQ49g
EWlSIpAbVTMuQ3ip6/I23FTphzB57No6weyW8/zdI18TdPm45l48HkdiHLPnxxLh
MmYRxcoDf7SjVjpMFRYz7eLSWrTIktbmWAK2SwZuNJjLVZlr1qDa+MALg0AobJFU
SJGWRm4jvlM3houYhCgIitp5pfMz3Zozt2hdCso321sJvXbh7FhyxhNu6aEYXxjR
67Es8u+uFsHcZdo7PQ+VDYHJduDuOwYgeKZGzNwIEeNnvWp9VYiQ5szecOkAsaPQ
Ox5mF75Y7Ju98hjs7dTUfm24dWF6wZl1vcDjj04nQnQ5JxNsYR/Ehfvq9DZplRn0
gOmclGtdtFVSUupD/st6DIUDrbY+uChLDpsq8/vh7gHJIursQITYgJQ5fWpPjPP6
KExWIHtGjStQkOW4jLVWg0rCKccH1ErglGKgruV1Nut6EUMrIKZA+RSR57XSbqkk
p2HefGSOWX8DvAmL0k3ps3WOdP9ywh0b+Nup5/0PrbkeGRLai99Av4SMAHWsERnA
OGaiPmVnpfO6Q/0SyATkYyaYrhbCoZqwuvDQrOdKcgccYSxyn8Buz8U9f6AE21Su
uI+lWdx/RFIyP7H/bIBVSHWDcyWrwBH+XfjSIglNyXY5laMyWssZsSBtgi3vFi27
UeWDhxEIp2rOElEESsmIEwEjfyXPdNq/bEjZrlNERWz0Tfb0hGA0rcYrApn7aWZb
APA8INTkHT0JoW7QBWKVtRKs/Kcu23E3bgvdKtyvsJnVQTzphS+l5CtLewkZgoiT
iu+/Tla0c/7AI0f4lo+c0a/zZdq6Nucm/FADZmEv5Ohq/gMjB+ZwYPC9Dk0BxvNW
q9dk2DxQlvfe3K4XRz6rLFMsnQF4muL9oCfq/SgS8B9DVDQpKn1xe8SZjDvhKGH8
M7G5pyIujFYvLp5CKaxln5tKu6MdfgstmBBwawVUEJFaNz/WuiTCzORLJ9+Sgfq4
ynT0mxLiZXIedOIQ7UCiz1czMM22lFkR8saBuj6Urp/aWvTC/DBQdGNQt63twaOp
czXMHV/0k1ogcfEgpP7cOWJt6ZlRp5Yb6YRvi5PJn+rLPtyw0jyeAtg8E4lf6Xez
G8TEvD1/PCQMypQ5IGAmr5qwYK41cvBB40UJ67ceA2tC7z624rel2K6Mi5xyTeqe
MRcO9dQpXz0EmaWBgzU3Rv6T04u/S5Sk3NZ8IHlf8sh5zgV32/tkVHxTK1J+0VMJ
mRR1zQOW3oZEj0VsFeBUdtWn6TQ3abdO+2wxRbHpmulufsvcYxwpzY5pHy7qwBPu
1V26L7NOyAXmi45ISPuWAsxrzlPlQhZJq0t5L/lunYDaIE8gAb+G180R6VzfspCi
UFa9/8Sjb75U5Z32bv361kWsXKNaectbdMpkGYUoHbUrCK5/iN4zALKjC9d0AR3U
nEvv3JnlGmoeeeDiXSIPN3GV3PLyiOsajxMVvzqzOeOYsSf50LzmAdz96Jj4sCPu
Mb+VnB98GA0PX1QtBVtWGKlqO/wv/Am2WxBxZhX5SBUL/EH9PSE/kvQS5hSsxAm8
Ynz3JaFUhqs5QmTh0O66mAnvsLf54oVaVxWBtZMUDPEpnd04t1SWrqkCuEj+MpjM
lEB1GFr92JCzttPu9TVQb7oJysspjQ2FnlUpBkFblN4mzuBsds58oYUIBINX8Td+
oZuV3jEEhgwWw7Bi/aZNincA6cVhrMQvYE1N3QERZo87hFSJidfLm9n3vdna7G+L
9wnUAEDOOG/n5uJKLz0ioffMgMUWM+WBxYDjImZKkr2OG8XFty+FADUwehW6qOHl
OdK6NYC45N4oydFHafLxUyiQbjdUzH7kRO4d/qmr4FhxCyMzdyZzJyBckkNKzZxy
4lhMICzLizNHmGS+8ITiuWI5Cp64CU1nhBxrR1497pQ8gHz1Z3Q7G2oXl7oWiDwO
L28eGdG9plstVVZix4WSSzWG0lIW0g3pPmALtncEbK/fwiY/65kBNLQUEP6iwwAr
AkOPtr39/CnX0/IUg6JA5BzXCEjuIPWF1Etdce3OD/CBFasU6QQD5ewknD2dzqmH
R0dmQKd1hump1qtoIERaEf/aC7JxW3bx82WPdQhsCc4ER0dUXZfCVYse+T4s7Otc
JXGV1xvGrfmW1KLe7pNKalo3D2vN8He00lOhJCkr/X4AK1HtUfIZyxaXZzIwOp+/
H7Xr96no8FwzYO8WCG0tos6S8SbzRXy6/SpBMJzhd6NInSkFwDfUvStkkXDLZVJs
7BRm7yJuPrMXpwEFBOgNeiNBK7YyXHCgVNBXplMWQiseuap+KeD9uDzY/tMKmL+V
yBGRxs20CNyhLlmsR8UFtlLq/h1oGRQekcUU0qDX1+YnHW5KXEIdNVO4M+HdsnP6
dWCzpNjbph3BU7mKOZOTGyoYyXoNjBaEyvjZf4+MYdX086U0siIDhUgimUAyQPCd
v/409GCYaf8DmgXT3oOHx0ysVZi8O1tKH7qi4FUO5HLVKEFUlk9cWM8x0lA3Z3CZ
coryh5IpW/OD3qhUMFVbtFUqwGtzmSXmfiLHc5JlR0IJRKt0ikYpJ4TrxAFNVRnC
CGRqTWWaPfNcF8tnKvjEuepXDoMLuYmuSxLAczh2QZKr8SgMon4eTLOmN/ZefRp0
0soV8oAz/Ap5Urdil0qndA/GXtN3wqT0yGuYfLoJYBmvCZnhApliE0DIAtDMdu8O
QX6sJJ0/pwiFpX6+bSDATt8wjrmtLIYkWaqW6+whljEMX/YfxPsxFKJ+jRpjtAzS
fHeM360vm0z01jGM9UjjQL1oJLrF4hqEVn309UHcvnq+wud7Bma6twpyDjHKuNh1
bz98z1mpWNMT1JEdQC1vxH9RHu+ealMt+oA14sT/S0/PbR1E0gGmRPCsMkwukWrw
3RtnovsWgq0a4jUhiYeonRe98bRgz2SuINY4hWSytozrkVATobS36m3R3fUxd8Uz
11WfLwYlqNm6f/gOKVMIq39g62hDWnT8mBn//7CLFeyj/Zct56J2NAadxcH/no2d
67pkDTTKspQ36ndES/Hb0O1+e49P8WZrfcQDt1u8XUW7wn5joyZF2UguYHtt+PsB
gofIedoZiuShQnylRnuLERlcKkV3zACrNjdMpIVPthiLTeDX0jE5WUBV2k5nVNJR
fDJO6YCyk/XhC2Bf4I0iVVwp8MzFFtklsx8I+ACVp7thK8N/APRpYvdyn/1xmNhn
K4sRYaZaWZYpj9KFnate4v6Msq4TLd4ubMQK70R+dLd0uuIj6P/sN9axlLUc1WJ0
jRlQ6p7ZPaO3w+wS7zCzlSrYcm6CreZsSL3mp4CCLQnFTdJx8wFv/Jr2TCub1KXB
ZgloRGixto+N08RC47kHsP3REIAbgA/ez/DPHXlurTDN/B0Z+2KMx958odrz8G1m
rSqQ/FkUWUQYfBA7kK2n8hQUmAF+yA+qKp5ILQ+ChQjx3nKrRDKI+JfvcBvFhROw
x8wApZZyMj0L+RilCW8cbWEJpR84rfkn7zFQF1eRVNnZMzPLYQnjT+i4vBJGtNFB
p2249tfIrIt/1LeQwf99/tkf/mZRc7Fumnc5MBD2aATihCnUUFxpK41IO4GcyPV7
Kvt1bYI+sB4rCigl5t2RX3/qoSG6cM+AGAolCyCZ98s/r87cdR/+S16jv8F1i+gJ
kjXCDh8Rh+X+39vfzgTVATmUL6PeITqvvoRwzez0MtrrCGFV160E2rk3LlYlIjIb
Ce6/c8w3jdnFSdhhVR46Fj7IpW2fVETVnHPzaH6jnb05YohaKp6ffWH44atQnDS5
oJBX3oLaD15/iXYIx9HCJ18Daq2hJ+MtB7jz+Jd7Yp52095UNqxvTa5hFAoJzkGx
hmKCnS/z4/BaDq9+eS/shubxPrQX+zZzWjDg7WGrRc4IFUQGVxVKcLw3PE7Vdp4t
0R2p7YWpBVJkIIWz4YFblUshMEIOZknlsIJAKCidWn+/Kg+cenipW4kKf8jtRhgL
AuyCxE7Jcan2+Orm57OGVa9ivbp4T9riS5JkTp/dB3IqYiXF/lJuCU7lB4dbZwfz
tCU/MYg3mGgwJKU07phwOcQ0vIKduMiQ/hUuhAFf8oDdDS2IZ5Urfr6+IosPOUsd
JkmdTuo7dEF6kPpQFFr5jDf/7tcAMljGdY/rJH2uogUhGQCMFvvCxHvHlLFaA42T
egiiCR2wNoISJPtchGYddvcyMrL3JwmKs5hjKsMGYpGgdzktm8QeQe7BCGSzSF0A
T6pkOt126DjaxRHEqJ78OOVLEALlDbBrPVWuMlyEbQjC0LwwWGeINtXou7zoxoMi
LkkXeeb6XHcdcfUjWQVW6hMyiBjYr+8RUCHBtpmPvmbJBeI3Xh332enjCKr8QeKj
JWtEGsU3SZVSINUpqSU6sYOFsWhWq0cCMFZDGVapI83ZXuYwYxyPYClXK5aPhk9a
gVSfvKr9T8ZA8MN9uuhsMMVyyvjDlH9auHWB4O6txXrORvNPEJXVshf1yvRHXt0V
Z13kGl0YKinPj+D2nqYSGw+ES5yYW/m4JoR2SkO3ylKGsoVIJMljk5JsyLnFd4xS
ts6eE37DoGbAJzV0btvtGv26R7ci94pbggc8S+42XfOsNcrjiUY3fLgnf+ms2D/b
Gfo6dIUIf9PWALgFznYPvVtf5SV7ElydMAqQCsf03wseqgtajyqIL3D1mZ5q9K0W
i9qoBxe7h/3gjW3NkLsPhdEUAfkFF+EAzQaXZgYnoDMfywumy1GeDdKG8KnpkMxL
FM952+zCDZG6BFgdSzad9Jt8GTT3xaZsT70f/8rIjzxkR1r1fkrJO7nHhRSffTx7
mSIallQm+xR2WckRso5cFSMI6kVahMLfZoDyaKbvtM78V1iatu85XHkAXPEEvoPu
4PdGICbJwGPZpkwPcxeacHzUCtJLdHr8e1JG4rv6nqzvZXWHtS924ZBGrx/nLZDS
LxRuKzetkvI36nu9V++MehL0+MrgHGclqNThpxFOdc4hhJKvph8WBW0Y1wF1kFqm
IbqYkXgJtsuY2lDjgkPCrnQnf403LuHokRDo7AP9yewTuK64VkZRMFmdEVzJjik0
SC7XgjbB0P+H1BaFKswAZadl2Ae6iiBd0yXQoSEdhkac5A5j/jilhH3s3spnJjF0
fKFNaluqqLqDgRCUs9HcEYBQ6QB2+XE93flRu6nMNkKQ5ihagCl9OH4h+oP3co5w
q3doED06BLoiHxbb6Q7MnY+OnPe9vkLKhCw3ts9bom04AZlvIX+wcvorkRUJmW2b
mLYWBlUDt02hcGWuPVjiDj2WqnLPr5ZgNlUZDugn/1mMop8RVS+JptE0UqiSMEyv
a2pMKYCBg1jj51vsOQqc97aLXvQeafcmpbCK0u635Ge4tpj7F1u2rMbzqX6P/6DC
dsZvKYQRIPjOMFHC9uEx7l6uxhExsVxz8EAP0COunqG52Vd4v8DKB1gKRmqPLbrz
Oflnt4vNf+rKpfd821trxfpUG1hsgzvEUrubMoXfa4MSMmyTBGVHgxw0OIgv0fAz
evJL1U5BLND4vhbKadNBOrFLoGLDoShg3dC18gYxIf33uFuFPzj7nVvFxFXeNPWl
NVvgaYbbcHmrjiq9CoCza2QmY3TRDASGANCLdBKj/XYdmwnwJimu/ExYJivxzRfv
OcRiFwP+TBXIIuxNaXEy0b+jxiHcXhySVXDJE/y9OXImTkAEVj8zppHf8YhTz8Ce
/ZxNF0YpEqCbrf7iPgeiR9aMeRptGwA3sUajrcJnKHnDWXL4bdhAIXbOCA+LcysM
4G+wUSULizj5LuV3e5bpxK9joHSU30Bl2pTsMnlV7CloBFVR3lZqJjmY/c+Ov6nu
ZFRTXtk7tKl76B47OKhWEkyfjQ0kOSI+RQAkQJKje0yDXiaUyiejIP8SpjPY/MyR
zOeal+KlPb/MvFDcDDOoOsvDoi5rkqtnKFBXH+7zy36TcS/bXj/GaHWwzYL7Ggb/
W6KZKPwu0D9LgwlBErNKSv9YfSHg5HTvOgNxYFVespIWeqN41yMrtNE6QSH0N4NI
1dy+XcVmWJzCy+ehszfmNghT9nLHvkhkg6DVHnmg+xUD7faosjDV050rclaEuE8p
rQ+KUc0e6dJvVlqprnlY6h8XbFH+YZCsQ/j2USVWnol0D4VIKt/OW3YnLVuCDDUi
6PVodLYydTzDIqKbQyiy4SknLVQhAUMh0BocidK4lptHKK1t+cAaTAMEh6fm6nUZ
nNJCvIJMzblT7bl7UuShIl92Sj9oYFUsbQET0kGh2SpaNRF3jjI1N6r4Vi8c1uaV
wE5PVT+qARoIEcdTJQrKRrVTPgeVOKJQ4ABamgqGan2g+3udnXqryb+Nmvo2zC6b
deoXlqD3haOSHJiA2DT4y5UR+FgssyTnhua7FMvHpXbc/JXYz410SRVrMPTDs/HU
ZExW54vCLxVEULeNfEy+AqTdlkJDg3hSLRpLQx80NtEfVHgSq7HjClsLiPKvEa14
utQ2NEAX1+MtR+pYXhXO4Y3vrYfaPkB6VEa8Cdft+SpOdysJEF4gC2e7BDuklpok
BA+EBu5ZqgJbRmmHm7o4tZNUYAw4adt9KMdYGNmtUCNw6A9AGCZKAbvi8ZtVq2nS
Vb+sd+mpHeyUUUalRKRsHVULmUFElRMwMgOuBHxJFwEIZgEBLUoFp2wBXxAe6Llx
pkbl5T3dUiI/Plr8vCGRYl2VNcBdctp7v/NBTplEEZhpRyRItRS8vpU6yhCuMfOG
ks3O2ONm8vK2N61Ax859357kvZi8Uf6nqPwjXLvolDTFj/s4OBYm2fnXuXhgvZC4
YgE89ffjys+fFeot2UFmNMZ5IGKGQZo8WRWIMUVz42m1R7iIvs3PI/4CBrjwtXp2
dcasoqgbGOFpHVI7rl9zzrQEKjIaF4nps69+9+lgkxwmqVFI5Ay33AFnipJodu/m
wRLYRxJfXSfoHki5hbvqOaR8OciBmDv6pm+8XnGDgjsgdfhWRKmVQ5dThBKJlzKK
YBT3tL+hUZ4h/Jik3Zq+8frd0N+o9FYmH9KXpLJ7TY1bAvaUCeUz62X3/QICIIQI
BKlEh+NUFB5YqLwjp6TZiNvti3lohRmcwX9Rh+fps630MhVPNaKj+hTB3t8Pdqbp
nd/hqj/SjNll3Kh4+OV7aMbL+ee3mMJaYianL/F8axtX+kE4ShKi1ft+LQJ0tQzc
iqlMeuDR/RrUfWQ4iGYxWh8mNT637ONfQLwTtOV4uoEAEQaedOeasRh4E116Vmfx
ulB+Y0bE7vhDknxYt4kcmUpyeCF0BxZy7E7EsWWKP5Dw5zEmnjSI6T0HRc1E5T4a
Vexsxj0XFyZDW1D3Qj5BBtlehulH49lB347wtcBRoDt+8pqtkLayrvyA7ZySCdJC
bwdAwyOsKYZrkCm27AGBR//qDs0QWJnv6VkNkBD5ZfCG7z5Z3xIOo4NZl9TH5BLA
qN8QjkG8iDh01NSgLArF6BZUrlGjbbbbwSG+b6zPoyQEgShexxtwyJhm/JCTvH84
3aC4HsjbO1GtfIdsvBdvH/UY0RDW1FJtXRcCioxIOu4G9eK3WY2YfTt61HNsCT9o
lnfqSFrdsZ1OdTPgJt0JDWtjiytdc5L6K9lhsfdy1N6AqM5HeBBzCyMKYM4+RsB3
ga0WO/vucTOm3laP1gN7tyVMdsHO6W65TcOKAK5AhzMsuSQHl0lgAINR1oLf37qH
qhFRDgG7gpcdX5Hli/LO6CsMOgVP4x844jaj2umE5PhV8tGLsVg0c/Zk6sVnOhp1
JaTUpqC5UIkNu8fogzrAAROFBjf70QUOKazi6h9bF+6U7uOmAFWM+zAqQZQQ1xAm
TrhKn5CRAjsoX5Otf+V+3heVa7y6LTSdq4IvBdFGq0LivZX4rPLkqstNSeeztqAJ
UH371nRliQJoUqmqafr1uYjK01uc1VdyGRlhCNKY8dj1lY8PyqpOVwhkYTj81i5L
D1Ycqthkc8CVmRTeBWHWyRO8OdrpdlPsqIGQYDdfKyyO2kCAENjKfQwhULKbzHaw
HMNJw0LIMzmhZPoJWPKZqtviiep6cEkjcg96PPxgGYPfPrjfjafQglpbdpj1b//E
0Nbh0epJKQCFOZDn3Z7zi5Gk7VTMqTPSv183FJ0MUAS9BOcUS3K43vE3TRLDe3W4
5g6NBhuu6iPmlM3d9/voYePwlXtLVy4OeotB+7I4WjS2L58TRR3Mjw9xfjoD7I/h
HHKR1wF49I5XZhiPw/UOtykdjkFKV2NemhjCikIF5N4MF67oCS/FeGoZ+FTaVJ7O
HoK1ymp7/JO7CNSKIHwFE99msl0DpAyIqvLzMSdPs0bpZrDH0FYZxGiCQKECe/CI
gEPjEcv/FFlJw1lgPTEvx3K1b+LSD6zOsbSrmeYVKRhAOe7yY4ykLXJ39sNbGntn
fzW+VTk/YSyTlgwLwk+AFMXpmmtNLly1+7YgETrNiy7abkRjoYPKhG3q8LA/uZgL
Uyck+wS1dA/OW96cBjvxVXGoKIiiD8FWCDP+lmVw68KVgK+kBQDwThk2peidpQI0
lm9WKesPP+kC+3h4AEzdzmucS5i+ZGrCEmsxVHpCUGx6iETCbiWouQVMz/Cbozfc
OpyVHXYQHmnjIgtQ1PqznTOHGGh4WYcGP4Ev3osOnsXO9WIhzfDludgkEkVTkx1P
M9xJ5JtnWpPYLU3HjWtBjm7hEZ+D8Nr9+Waqa3DC4INDAia1L2/0cBaBSPcWTYQa
N4cfCSP190z4QYNT8J+V5nm9eeFBBL6ltHX9VTP5P6dNclSnYvrz/emEolyk+H+I
96ILdEnh5RvBF1ZOQcNw69atPyDjxHBUtSu4m9gxJ01rSmRcbGsg90b/2XqdE6UI
EMPC7hbv0d3U+2l72YAS9gT8w6/FlrrTu+3tiVe3/eyQ1Auat925PcgE9l21rXLg
T67ME79E9CCnxLaMM5YJsnVCJ15SNMHo/gMQJtqvAMWHNUU++tVTaVc+Q7NWv/P8
4UjdpqrZQydq/PsCM2N57QQC+f0ePqRITVrJSTgzYPyBWqQ7uFCjXHuGuyxm1yF7
3ybQWzNRweRSd2nWGvqLUxsQd8/Yg8phw4m+sDDqOhLaxotnH6398LQsdRNG/DqS
LgWIA1XHp737MU/oLH/vPch41fARTcUgfVP+P9Rzf4LL8pE3cQAr3aENfMVHCOJ6
9RsqvdoFgpiCZOf00qOutJkdNmealObnnypLP2bC5M4h666BreicmmYXPQoJ6AlL
Capr6xmYMzS92Cz9fSu5Sn3Cf78TrhDRPeDFuOuV5KRsCWWWO/JKDSpdnrIYFtO+
vJpTRgqzjHYTbQNAjRpGJumDmXkHrOLZbK90GPpaD15PN05wAroAlmYuzw/4s90C
r0N5qwqpIdmqlm3zsW2A70sayY8e6qyiHy5h/6uPfMqjMTTHnJYZlZjpCX0pCBF6
JopGGalwuznCXbGz9339HQgcIkXSF9LP0SRB718Ljzhs4qRkMQGL/OLvso4eeUIs
oPob6YKsUkw/uP6NZys4tcBTI6uaGD7bVDy6AQvClwrLOLSEVeN1xQ9qqilHagF5
9Jp0yE9S4RBTGTiyvKkjthwwXsckrg/rX1rLFncpOrtYVcurNK+fUCR8T/HMbHck
9Ts97oleGsvfYFMDfZaNGowSWasWuz8Krj3rC41gtbr3jonujImsSylsv8qZQskc
SSGbSdNLJaOibNuvJPx/nbNoB9p7C0A7lQqQpSB9mK6YUy5V4RqanpuAJm37GN9O
QhUunPl+QaZGNTUz+eRMUjksV7Cq2YEiCv1FQfhF8H9qPRG4/H3zM5xqmVx8092Y
jABpGN+x4P0LUyWhSqZPXhdTUO4e8n3qVCKv0Sl99Rep1SUr9rtxWanOIAJo3H3O
deIQerPx9yVg52M4H1liekv01TDzih9FZvDwyflCZwBizfCue2AWkRHVhVPG25Ka
vf827F+Wi5SXyzeDCQEXxaII5oNODo5U57IduVr3AUWRQm2DtAtEcqDF8GQ6994c
nonHxu/6vUGjGhaMqB+o7mE9UcBLIvahFS1BQLcDYvg8VrmXM7GNaI8+46USpEHc
nBUNWZLyqKQzn2eKc1oArLBWmirbxZQNphNJDu/VfucLyIKwTchZ176xevOTSE4Q
1svbCjo0cbWpZVL7A8teBpGkeNM+80e+YXTORUnOAABbyGrx7Tw4GkSzKb31NUJm
fwkB7+tAfCxGYYAIUHO1Lt5POSeqcdsFDv8Y3mtOi8dYpCJ0qLvhpeBMPsda16dM
EWdk1bT5Td6KenRTxemM/au9cuobtbM8j5Rv/sNo+ixuO/E0X9elO3Htxs4T05f9
JOXb7LKnOX7WJ6MPpme7VHi8D7T+YXfNNlXJlqiUxI4P970IcpzZiXWp6I2727Op
wxg9zSY+t6ZDdhC9IVzFBAbC7d1j6VrHrUw96LOUeVVp1HrKk4Sk8GwMyXg0BKB6
W72TNBP3+Kc58xTOAHIX12zqKYVKizY0SbEAmAo99U3+8BnUbPyjTB4sWQgdsvbC
+xGCuFPpCG1v78PPTe/Y+TZUkShQNVFuwERMa60vizgI3bhvjjJoWwgkotlswAIt
Y+zup9yvWy6TxGj27PIbZJoAWggHU1UFM3yNvMcKKUCHAAH50AaWAF3l+vtYcJQX
S0rfj/M49AHBwYEKd7loOS7MVCfQVuTVrxSUWBRoQnFye1TbJth2Jy/CzotZQk5S
NbNj67suOaYea7gGYoj/HNLMnaBEg14i3qbaMqs/0DuFNxHNJwS7p0xrTAyF17ni
04h7bmeTKNt2FAoEBYj8pz+4BKFl33YRGoQzskpB9Vr3dhTRT39RYAHW0lxNY4it
8FdYQp+kjQiIedVKzJoXq937+TPFItE/f9SjDtPjZ5/X3l5W+cGctjzCKy0RYbXy
l0P5j0y2ONZnnJQT3JVruPBwSFrtOzLX2eTRVeGeLoOxmBTNrNQ6f6TuzvlMR7Ti
bBkHOvKF/PuWhopFggtJ8bsuK6yW9bW6OohJFcfp+O1ri6qgZTvInnVfjc2+3DiC
a2Yn9k3I+LDJ6Feltd0FVsIBiZLr67IV1Igo0NrT6I9AxTWykLQaXzgzXizdchHn
eOpr+4mosJf7rcr+Lsc6+bSXgnyet/6cDzDy+VFWzsF1e7a8HiqfKXf6aiEYQYnX
bHakEU0gS0Ino1L2N+0SAfP5HlnTKIUE18hTEZazP1NxtVgYWPOAR++qU93KkgZ1
hlh54hJKmcCtynip7qpdo4kO/HIe3x+njRMhUDYXOWoKwP0v67qfLAw+KeNsD2mG
HbI4shUCFrxaBL55hQ7wwFUBcCmi0nieZuTwtLAmvwxR3LA8k9s9TajRqmy/HWCY
DyhCaG5QhvV2Rbzjpy4nEJQ6mgzWuxtznHK39EE8cNa6CR3h+2ZBzT3UykyDTOxp
uKJLF6vNXA87aF5lytwdIM18DR5D/vYNhL2/g16MIM353+kcvL+wXzZA2cU5kbb2
8CGI3ahBW8smmqTrmy5Br2YU1igaqtFy+TgF4H4GhI3emhG2vIz6iIayTae3bd61
FoWkQuHeFGIy6znsmLfRtyur5BQ97lRYqEuoCY6I0eJnc4G7T9fzRQiQp0dppq3w
1EmZ330BxtnDxMdhOlAqdMQUqr4S2sUK13GgIKywqu7mVBtDMvclQm/XiAecZTz4
4up6k9OsOKBZA9NmfsNPkXu/Uy4A6oShnd47fgslYa9ZAA/1d+OjFeIYtE2kd1eM
7a3csa43m9oTI6Dvi3m90aJqw50huLub2B2JuEfcoqOMStix7qO4aUrb3Zqomu6L
IJ/hC1RtoBCO/o7BW0w8Xch70ktIFRG4+N1xZUvp3qzK+WKWkG33i1+TzcXUbt9I
pVb8VVZp1z8K+xf/DtetnjFkEZhchYYj+7l9oWdVScDo2TnXh4W/tU5OBCap4qAT
dTl93QMEJ1Y1hV9EaDVIFTanSfxV1lRzGU5xyeR7fhqIeLTUxOBmt9k6iv1m2TSg
0qEYue3K6N0hGoFbv0i32jrKKfscZbsP4CXE4FfDRXeBiNm09TZ1E02DP8v3xQTY
vQPrYu7c0cQl9pfC7ndq8sVfGlzS5bB1/8LFtr6lFAxJ1S95kWHu3F/W+cLHuo4b
YeERMglSmTBP2F6MPHoQw+UrXCS1jNa+x9YHbLqEztbnXTtFVPiHG9y0+pyCYdZg
08ZM/SBM2wWY0Gl05TuXTNCtZGQzXjW/pLP4rSDGUwCuY6vI0MSTyPPybYfyZeSt
3e69igQfg2WTy8vADtyTSW962HKEzcPsI+lpRWunaj4vXwo/Uh8RYS/blVA8rAoR
71q8Ov2J1fGTJTBCh9jo39dk87NYCbH6rGl/jsSoHXtZTxW4pKVuAG/p5yUVM1bx
H/Km/ClEQ87R9cUFqun+YufIEjhj39zPR8kFSjozNhWe3cYvzKwcEKUQzZzpRnsZ
UyJ8qjU8Gmhs1SiZy8izBceneFyQK+0mRsnDFBBU3r8PKje7ozW/JOxWyeARP9Y9
NE9Vu2SPlfZ0j5ILBKbK7tyulmdfgz+hkUlNDUtOXPdYTSwb6nXqQSYKH9YhAPkZ
RXzxwTOWG4mmWyRbPUUHLElkXbg6+vX01uu+5VyRzJrzaxmQJedpem/EWbMYsR48
0/JbMU9PJX4x5L1BN9zBqjASOQ1ESmfw+9iHXLNJC+5hwCB9ZcAra9UiYtDKsTyd
7xCF/867tEZs0mUQ/U6on/Yu1nb5uV4t2A0QMFMrYu+A72M0WXGc7CQ38Lzs8VS1
CfvbNTofpfPcQ4BTLoo8kalhvkxYrOBfZ6sa0YEz+vu/5YNpvmQLnYO0uB2nJxVO
93pr5JKnA9dGhw770esP0Alb4+BaGoIhrapCcOyDP+ne8fpqswlmihznUGWZ0WEH
+Zqlqv8EAQjqM5epJHUqslYU9GNxI3m0vgLDTzc/drxQe+80lqcnxgWl9WgIFTvy
P1U93hjRAgFOn+6/+qjPnfxhmRCPuBk5B5D2HtMpq7tNY1Jar5aQdMv2bkM1IyCx
301BUc2qFqBLh3sNNNxHs7T1e2voY1p+E4Umv6CuUkLhSV2LNbIpdhk6a2t4Zq5w
GXMKOdJ/7NJz7XjVvy9p12D809TRE8Rax+mp6rAxxQZMpJ+58CgM+HrkUC+Rr1aO
sd8w/acoh8O1gYQbuNmCfdwNKFuyVOa/fVErW4PWFCtQfs8sfssNLCURB5J56X58
64G5DSV1lXanRcDrJgvk2c1ctLLgXyV5um29tBDmp3EBZZbItsBQ8EFiMbZMoXzT
jvk/2U/787ahBwcN1v4Smxl8mNrx7DmGP/RUDOtkSEVLPynKr138r6lJ8hsuXZot
ZbPQzscyGmR6D0EXJK+6FtgzZi4hdmMDKA6EwJhGlUheezEVPYMdU6yfuux6ZrWL
lJHAKsh0qkK88LG5jAit8xX2rBDm91OEctgmBkFLZqo0SqecvhUuMbxvXQziw5th
SMGC8WdyNvqNjGO5ns984HBm+A2lENpUH87Hr9WkStYWUr3F+qKicim5wt4MUG8G
W5HiXFTPhfpZ8NLiGML2NqSRUAx0+ALDVuCflnPQEy4FLcCX6eLdSxrxB86uRprq
eWXCgsvTX7vJstlFNysaYvLEM0NudN17jXRsnpTwduph1h4GDAtncVivhYftENsx
zRFPBsA4eJu7un4eInuelQCJljXC+LXU+AkkbvilIg1/6jWpwqD+ncOcBt1n4S46
aTwI6OstAwAK0MhuO05RBw1j3pCFz2WAk832QFei/k/Rl2b8iY7YL+/bBl4lLv53
+39jwDXS5dlQZ484XnWq4ZSUl1kztARrkDcDSnzQK8F7lcCIn0nomdORHZmFUecM
RD09o5L4u6t+7VTryLsnVg3hkG7QmrDrr+gLeYXTirILzwFwBKS2Jc7pCOLsheK0
sNRonS6ZNESgbPFDi6mgkpTKamWfNWgz73JmF80DJrUaS9/q+6mSHzX001RCez5L
ILTinUjDofOlphJdLCWb7EkKyEmMiF2ZE0u0DM1tc6MB21t94kAcjgRosrGaIoH2
n/qeowZTa0HTnxEXrC1rK3S/muwtJ1wbAq/xEPt3UyMx0P+FwTDdJ5Dmf1CEwD36
t7lyo7ESdysO5MDBWw9445rZGHlxc8Uce77cBrD6MLWvG0w3zy2BthH9J9svr0oZ
7yemHD22FaFmBJ3u6FjMbs7Yfeeip28AJF7jTXJxHcG7Fr/BLxJB9NeB+PYyP/RW
ThPv8cODwRR2/7ydl8ayP8ISD0JPmSo7N5V/62ALhN5+OYY6EAYVZwlgIkhT51jl
2GyFPGat058sl9bHwpTA++0qmGBj+DiXqjedfwI/tcdRPl8bRnuIFIFY4CPKFM87
pNzvyGIAQIkXDN4JLQ4WLlYPnW/RsgE/KF7vsTJOL5fqckQ+CSXj5YlI7WPNAsNR
0ZyycYSUU53ZIFNZra9UmkjlbLB/+FTpzJUMcBa2XJkLYjFwP56VtlkpguwQS3RH
Hsart9MDxmdEh4b5ppVWNp/+yyacJ3rUR5Ae6xYG/nxNwC4hWwNpy6ocdt5H8vq1
q9GNKqrKMM5f7gkUIuABEVQujdGYw2/Nu7XGABEPtpguEpsEfqQEkSOdNPvb5pZn
91YQPN0kL7igcZjqTQuAE8XwkeDTr46DkCP2na+Je8atFm5DL00uT9T17lFCdKEM
qx2dZihh6Z/b+agUQX1HFFY6xrEQFMr67CzGX38590pyanNwkoNH3tuGdOO//r30
aLLNJ9BMjMTyHzWEJMySgWL4Kkdc6BTITnTbyc+LWuBtfjLAjuXToXaI5U+ZSrFJ
7FcUdT8eA56AApGuyXlEiR016pwRlpDgx/gcZ5k76O6POLGBScOOclTzR4BIrsoa
OoppBhy3+cFZBwUcCupI2zsM8vP6DfpyNt+fDfkQyor2ZFrxYMyCAZ1hXNfo8tdd
zAfhOtLBbWLEpZxthT1l5iQhv3usN1POYThm2ZEIWJimo41cYvy23me/CfNb86FA
Dy+LK+1jDJ7AaOKKRyRAeAa2iDnQwE/b3/Hz8Zn0z2iJpOUnA0xaBnmpb3iHSnul
wr9PHYC/HeGVeqTurSdGgii7wXNtJQzddnR82swIFtK7HzK7O2AisXNjtjAN4TSX
rPjV5S4n4khxzAMIoN4RbbComvnwPYJPzZvyg48EwOPBtZ+Uk5Sb/dTvm7HwY2X+
JIo34T7zI2PnPJ24QeAHwXCwsryV2mB65nAJw+Z0V+PBAhuwm7p7Rjx+k55dJRe9
paMsURKMCgbmBo33igMCW0mp139Mx+XWyrTei9Jj2S89/cUsblW9AXD6e+0yejiK
6Ueng2roeIYJzeZ4fMWUCssCpZzlXPw7X9pQFKPkT6X9pSM2I+nHszmLl665aOck
49YmLL7JQl4Hr31zpXZMvL4vmt5IKNwvpaJJtRmvcgxTyh1XQ1DlmoOvIt2g5izv
WE50BS18XHbnIdaOC5q69S6PpYsMNhnsUS80qD4YJ04EQJJC36cYUGV+kA8Bh0cv
7YCIwdG+bGbZ+psd/RmMXi5YN9y6yKbpp/bZuZSM5/Cum+nbeuR/kb4ZdH2juqmQ
QiYyFdMXpU+tmvzyV6vcnnyE2enGlA5Tqy6ssCGzQDkDNN5WLlhOsm/J6NDeoQ4b
sOU69sc2OovqAzTLC2TkKeXemEUC+tAQjS1qxCPcTv5K0Tp+rCQShNO9gaySzUet
7qJ+Pr8JYV4kqyIL2NFpkW/0vOutLRxBzTLQ/Ehs2C5TSgJfM1zUsdmTUWXQBLEU
QoUmxSRvlpacz/WswW20Rg+JZJp+9H18LHRInRPl16NBirPdIw5ejaWJhOJ5UP44
rrrG7FjYjIDCry+IQOb/dm0YdXaSc36BUgDoLtVmrW8QaMFms1IuS5QbXCgxKbdg
YHtRDvSjIjkpqrAICTIjFW7+RfZe10t96hKrKcTaoFZ0/ZCT8lxwe4GjRBnrdAyh
QgHWRvS84/2VVxSpKQgxyZpHS3P+wrH5BfMhog0YAsm6rjfl1FMhUwwhJrhGVcEd
X1fOmnrNNngCy64LQF9F5rGUJozlgK09+xQ+yKkDs6FnLmhcgsPT5wKckYMeYMJd
FYR45cLIfn1W98nojs5wgk4+cZPt8e7ZTwG1fnHr3TWll5izg5518oKeLvI9R01b
ETOLbwMh3wPCtDXE1qwhnUA+NSO4unRhRC5VKiCcc9jyMLgRCIp1vPfShBrv01MQ
ekyferwhZsiG5N8UjJlQnpTUMQTPB54zsSg1B1buWPGCmgxhTs+koJByMHE6GcPj
lBBdFpshyW3hFb132Iyq2VpbwaoyBKi4w/9IDDMz5slbsXbcxEZBni1MQ15Bia1c
kdmokrVLDCMXzs4BpuugAxOR5/z81+dlVNgoc/qZIfPH5Frn8+F5Qrc/v0W0jfu4
u6ecnV6lHtYOVQhcEaRS3jgGoAcwPbFWiu19Utiu1NE2pDJY0y28wJm8t479B3+t
l5FCewwHQnf4EheE/uSJ1+8yovfkoP5H/rbZcthCbfzEpuW3jggKOI8VTCp1ktRW
S8n/s+fHkh1G+hWjx74nUG3qUGDjt3ZGpGs+op9ehqFLGRkcFeQ/MSUcAFroZKKf
kEyaYVRZXhyv8GzNu2h7wIm1c25tSOodi1j2q6v3piUP3FMTbVENZNPl6cWV/xeo
UyQyBC4BOCYiQH0JbY0TyPrq/1YlZLnRkbbH23CTC5rw7TX45Fo1vs+yK0FD0mRg
S0tIscLPulXNh1MpYZ0fMzwvJpp/Z9cjqcHmN/Zso/LBK5B9zq3OTMQnBxfx4Yc0
h5ga4/sWmzWCpLeR/aFDOAkJHDGTylZsfIYnfknZryy2U0mU/U+knSBeAfUb1U4d
9TG6+6Gun3mOPcsYN7TKvFp3St9JxN7xrRB9IgcYf5LmyYjt9HqPeUAtm1qWOVzj
CQEQrzPPgGCzVB8clJylIwfFo3V87veC0n7iq32aH2gJkN6NDSXmwGQuEjd0bg6t
pieEjMswCzEOfKdpcL9xsClKgMq3F/Bna1PFXR1ttIqWp5uIwO4qTdOGl+FnYLsY
/nS5J+XtfcdmfGQwd7muETwMqpfQmYvmIMkmxcNDi/JEPth0O544fCs1RsXPkLDR
PP9wmOy2EDLXslAeCop4if72lHli1VF9pQoRCgqCZH5MJKFQYneoIU7dP9M8NhPo
V2S7J0fF/iyQEU0E22nqnijB2AKzoo1FJVYKLzMXBoB1TCLRgUNr1Fpx9GHninsL
p1l60fN61DMYnnjGaz1LCdIjmwNXpr9ZPRKNtW+Yn6eWS8w1Prziq1tL0KuLBf+R
Mwwea58sV0NrHyjbFJzAnBtsk9mbAja/OqdatCwDjgAQS8nePI68sIeXyRgFtI2c
I+TieYbWqW1XzkxkbxeZ0gZKWv4QDlRYp4MWK3gcCfGU8ZDsjxnHEc2KoEsnHXff
+PaTG7pwB8Men89GOFpyY/Duup5wFAmpbgANCorTdfjHT+Zb1TZBVDXMkRwlWP5O
xfuQfwgthinhz1XAWAKheEQM/ylTSdPz93aNSCk/7LNHjeTbQfgrpw6fLjoIIMpS
UappdFSZT9XsuvJSBYQml1C7wi3mhF0bP1f5hP72N0ONJTTQoWAycdqiakeRprxD
+hPgUfOX2i6JC6tAjLmQaQCwCadckTONr6Vj0gwc06VZsbCOmCiB8YIpAfJi9Ijm
/qfElRuGyP17NoSfOyDL3KJztf2i0YRyNMm6mbQhiJFeA9UL18uBhSbiMEHKDzNJ
bDwsSyHFIqjsGxFx4mULXKwpWoloTham+XAUXedj2OtlfxAaNqINPIdTsooFhtuG
prxGGT5pR4MFagifloYVsWckD4GtrbyKjg+8C3PEqf/QY/fdkAn6Zp1G4B+00t+7
Kn+PisVYKsbMXlOCLqQDSVbNkvbVD4NCN0blCh3cebdG5KnyottKoKW6Mrz8f/Tm
qU2ZHEnytMmSyHNW0w+R69ganThaNwP2Lg7qSS+3q1ZOFxQQDMuCZ/YFBssiRH7V
BTllQ3DH9Xs02Skp0PER2cf5oKE7xtxjV6l0o+OavUpJM4sNb8gf3XANO2f+ufBV
wRv/8B+39a1NgfKJ2K3oDCgtqY7awEwN+TC1mQMy9+is5wGgYtpoiFX1lW+JkP6z
L1fpr16UBe4/yjDqlck/fnncCAS5PFsxqGbx23hqGWiPma7EWf1LqVA1XXZ0iFLN
mUGdALO28LT1Ga53AHitOgjJ7Zs2mSSKqc6yHnmrw8JF6ujoL6WMlrvzQTsUDPl2
tNubP7Pwu5lHg7sn8KuvElchBGk6vpdu4fNsKttx8rujOQCwukJ6FuY8YXV0bHnR
eJW2bczl4ECXWLmHxa2AhkGsy/2vfVxGpg+fhcy6ruDthgtifqJzm6nbSAQoT9XG
EFPVp+ujzCQxjb/vfYlJoKUwKi2GHUKlYgl9QfK6Zmq3R2RvcGD1UX23UtYzzGA8
7eQTvVq1iDwbHnN6jeQ1CbiomsvzN3ZunsmHdCVVLtjWkSunNv288iDStQmp6t/u
HDLZFb9wzLwYkHb//d4YWOsGyr58zCWB4Lf/1k1A6kz/B3PZiW3PhIJd8Ehvv6Ns
4gCXfN+6Y9L/Qvc1iPdxbmeeZbvXRmtXG4kMgj7a8KnMJBy3PJQHZlH3s/yGu2/V
x5I9Z1bD5H+G3nxOi2z6CXZHXUm+1IJpj9dMPJJ1EnL4OxaffMKb+FVXDLqV+Kz2
iW3ptGdH3g4531z2MdBEFriR8oqPB2nnoVSB0+XtiF6fbT/Ax04L3OGl0PPPCLEf
c8nFp/ZiLnIjdtVNRFqX6Q8qiueQVt+9kbkHSzGW82jz2VZkhYkkCOyK/qLbOs+d
AmBHk3TeIVqvhmrgyiquME+jXYKpj2wRBfQn/ZyfjkdNgyM+ZJrp/MP98rdVhUCk
1qW0HO50lXbfxr6gsehiBThwmSHjdNS01bpnRlQkpbym9DbOlQNGppQClRiz/R09
fmQdTUDy9upjhQDRYpACVbtMMxcImDYL9P9i8Z3j2uGgrBe5w86veBHCzTywrl8F
0VzrcTHvQaMwue+2ZbaYANRX9CQi09SxU4HRLqm4aML2u7ksGjMQPVqUtIZMWg+B
iQO2CxXAwtaOThzEo+t3XXITlakOS5qOaB81X1KTtQDHPWUWsyrNAmgSnoxK3Ocz
hS68gNMGxlnmD3VTqaJCN+AGa43H/pRY9dJvL8+31EqwIf4zMHQD40eeY19MC6nu
KrrzpG0/9vRsAkbBRUaPphwV9FtubqNlVKrLu+3GL/7mjQhEy28/0cy2Q//vuEmU
55ZBYjKOcE1HJSOlMPU3rNS2FvSBh/mqO04l7Bkp1ynk04v7IBcdZC5So2Hohwma
zY7Q8Zrh+fXVmuy+o+TJNJHlJqlYvTI78Ze7GUZvRusWjQvG4OBRex4KXp2jS7bn
cCLuGefoeSiGPvo04rSRbVWpK8ceIKerN3VxfS+h15LDZSAfw2IO9X8uf/ki1LrW
ZYhQYKBLfZ+rQu/zaAysyUFKtzRbYs5ziT11dAiTkkfId7yGvlnzTobGiVBYgAJP
OR9zd3hVfQ57sZ083q0jfEKKsEmwdhl4guiod70MnOsLn0z4GLfi+052NAYTrvMf
461N3fo/gqIKvRdppKMeVavBgnMoAzTUgWrZrS/scjRV9gL4qqfNnaIjP/xm5PMv
HiX+aDLKSskIwldKpX61KoTgv8dup868vXMRyt1PjVQhASSb0EPNb7wtSv1GEV9j
TKAIBnEFyWIhaZtHQyIH5fB2TJvzDNoSIfQb7AlUvd7A9OcAuUyOF5Hu/LP8BLAg
W4bH9hIeEhHyl37jgwKDp0lfHietF13kd5AZm8Q9odbZdqyJ8x9bcMXMi+jgCvsp
GQxPzRtLxAxln5mS4E8AA3fiVQLlXni0U5MBVJqGmxyLc4YAGheDy53R7y8iOZIY
Uhz9vbsGCEygAmqUyENlO/A4skwxdodTJPkTGZiYytAqrN41mgGn5/vnYI/PFvV/
Pkc7nUdyRXnHv3BIh+KAt43/N+9klQddgVYltzbei4g9t9LnGsXgNCJVVWHGF2Rg
6VGHnN+519YcogLdAbh3K1jS7Cwr6h65J35twhvIMv5FOjYiIZjxExY/Ag1sxweg
ZZok3Ix9Tnd5hhchcC6P4SejAxJupNAjDjnlc1jmSH0kfyTWo+sY0e4KLtE4NTbC
P9+fj9Mp725NrpUsNj55ZZ5t0HtAgo5eyvdaSqFNYwhkoNAGNBgIWKOaMBUZclE+
GA6pQIZ3Iv2GAuGb7zJZHnQtd5fi15SGJwlfRtU4PJNMr2sLpqWZ1K8DwIhtc4lB
gHjv6TBx6FekY/IW8IHFaiZv/MU9bQy7wBf4J9jjr4OoH5TGIMsO2GKG20fDpgdn
nzOMj4MqUCnvg4y+0zgebNGo9D207e9VmOOWUcpeTc6MRHjXv3rHPz9OYc8WCp6V
jC3IaaeecQOCKbOVUsEApaG8xiDePRMnuEBlVkEgcxhvKKEBau2AGvN7QpvuksDL
cwXGkdN/qp2VZG9mi/jIDGtoVfCmB0nux/2M1o/lgQEsIOYYk7xLZpTLfoj4APR2
i5xHRkhO27BoMLklsuNbmZBWFbFbxU22W4J15e4qhnMy2PVvNP1ERJAYFGMeTpMG
euOPFP4xndBJfLmKGcKUAykTXiC/2B3urnedtSuONgHE7YZ8oaJOCJDu0jQSKJ8R
fIfAf2YbPiapes+MAt4p/DCeLhAOiFP+3WarvY+ZEnfT2MX9pvVIxHuJS/4vx3t2
uh66KZFkqFzpg9S5cdHe05L1Cj1Kd68TVhxOOpzcPewwDCIBptHVaGu2znFDUHMx
D8k4tA5M4w0rfojixH/KXrzR01UkzW0IeRGrsZm2BpRBYTcw7q7GrdRpL7qbMwTM
30AN2d2Qjs3oxcBBWz4pHOXU8i6dPajua89xc0aM85Ep6N6XtcuxAEHD31gROsBJ
Er4ajMAUM+P9cmrim7pu9gVqdZZwYcCzFAbr0DIB1PI+1t1qk8SfDHHPVkJj2H2y
SJ1q6W4DSZFlxWMP0kwDqj2ved+AzZDquTXLRm/ZNUU5QcJv9u4ThZD7daR6+fkV
2Bpf7EROZlSkeh7GD+TyAUEavN2qv6eV82Nt1tMAnjpfRoufcjDmisOaBLePhLn3
bNl/OAShwmuxOr8xV+Y4b899jAwcbFryNSBx1cdIgI36HRznWZDI4LcDKrRqIVLr
J1f+btenuraQAwisF0DZgX2Cf/YDVpNQzD9Ew9dlBaC/l+8FLIruMXlF6J0AYqNL
/ioWXdS6bQb7zgz7XQdU6NhRXMFITfCm0BWux4ZZi8R1HUwfVs1aNlys8RQaATa2
1j1jjR4ltXompfi64tvRRHxGlutuheKLF+VMqnNgv+0i377Q/+STwOCdYdBNZk2S
ifcc8ipghpW5bzI4MfVKOtf4UMqDXRetqBqcn/NhdAIZL8EWqCwGwHRAlhq+y3fG
q9DqdxW+AGmADLqxRF9xfLhQXqtKS+uEJrYW5oQPECHtUW52bJVBLSqnQhR7BQoC
ACsYBCUKDWHZL1X/e3AH0lhbPdJeyHKtt8zBLkbV+vIRchiBDhWDXLD74PoB7eW1
6t+IlV0IV88wfcUpDvVPkzwNyriGk8OW487wKEX+KsruxbNzU3//gJRGpn4H3y8G
AsKfkDW8Zi8B6OVj5fFtFspE6zscnAllSpjLLvvKVFHxkdradEU9K3MMc8J0AAQG
UlAHTcGLPEeLxnY7N7of7W2THqnN2qVXHuzSQB/WH4+M0Grm2zS9Gn+Mv5AvouGq
uZ5EGln1QbYs1Sqsh69pRPOFaV5BOUzqzPns7uD0nLP5r2cdj0wFXgfIrPBK66pj
OGhDyRXP2b86Ub76sCcVeWm3xANpCr//f64vqfxQnA/RnvARgo/5dYXwl016KVlV
LUjWBQMKqkNVMwO9pc+xOrUb3y3obkHuTHuTZugDghzPfqWJZcMVIUDaSdwZjZcy
aDffuGoA0P6WXF/KWlqOg+tMdZQD7VN2S29bqZub1MlimeGejHo5ij0o7j93XcX8
E1JfGEXgVVFoUKKt2QpSCQ/6Wkz78OubcXSRzJExWIZLbRJKyYPDWKLhvnBkSSii
pvZqDp3Tj7JVETh+RGYeO622Hnk2KC+Cbt4GB4Sc02rKsppLkWXhoiKuesp2KM62
aoB0xmR0BdPc4X+Rr70atOZBgweu8Gu/q0XbnSq380sicFKO0vSPsDtn17TUw+N0
KANmBWyLFzzd1CvDkreZVkrW3Hli8NOvvUdxCf7RdHBdnphIdqTTAaF4/DrXJ8o4
J0H/bSjP/MOZWcEB9YBsvkxLfEDOEj5RdeGYsVZeN1c6UKJS1oRTbYg0bPQ6OqM3
rLX2u3bKnQ8keSWcxBDns8qsSdkAFWtUNta1vwo54VqOuYexEPE3sMqAz9Y+qvLR
MJYLzxaieRLrTHUxY7AlMu7whVqRruNENGn3xuNiatKNi5MCO7YWGCJik05GGr6C
hI5utLApvKQXTH1EA3wQujwWwjaJ/tF6SOILnka5640njKl9itBh8g7LlEy0aQB5
fpLd1+dlR1SuT2OL51LeMb2Qz0hkCgOykbh6Yl4xMzLrETCRnCHqAx64CED4V+CY
DQXfmAHMeUtC9yuLbPOoKtrAz/d1PCLKYCC6Sqpdji9ZXvTrjb0fyoNTeLq6OKhr
/y00kGvTZcAhY9xt3NOrsr6cfVdbc/sQiyNu3qssUU5RoBllEXJdfuSk1cOZv8h3
7IwFi5Pqp3FjPMt9K4QzcF5yKKAHcyK2OmbcOfUgFjpLGHff5rHGqKhwrquYe+uF
JBDGJKu2Rukyff3BwhxYBWFqG7SNCUX+ZkrnRfovtE7QuOy/0bPquR6XFcdj6OLM
Q4lAuG5+E8xQQRNQ4+S1kHRWTBO6y2yZ6evMSzoJ3bmyJy2/GM3ngjrYOfkB9NSh
qwMMdTsaErJB3musIlZLL+AkxKjTej7dUbac8BrBrVb2CO5MRnATpfgsdBQMmy0V
bT69t/GBDslXsO2Lh9AjYTYavdkuyCTu+mUhs/I1dhGk6yOf0H2LsoldZSL5zEyW
9FIUciQTl9Dz57KUw9FhG8mxIBGyXVIQwKu5d6w3jAmJ0alEaADQ1/9A0uZmXmEc
DLLNUOhUGVBhmZL9wLKXWIgZKE6rLpQIqPjAdlGdK3jCIEoBOeopqL35WyhB+zzz
H1genxcz+nlhAEf1FTpz92P8fFgfgOzMqxPJ1K+71K2PdEQwn6agdlsp4tPwTbaM
bhf9+Gq4860WqV3qX2m6IMcgvT9nTP5T6s0S2Kq9+9r824wW0TyjQ/3z1GWL3zZE
p77xVKc34JX5Vp5TElEk2qErB2pKfMbnTtIOsyOmD5Okyf7R6EUCqpiBp/TaHfj6
fK85pMTNoO1F/LGB+QRVD15Ve9XAdUZGPBd62li7I34WbWksEdb64wuCg298VDr8
PIZtUkmCCHuGEY+xaTKfyapfBhEjIEiHhq09GIVKFuWxaH0B+7jdilmZVswhTX9v
Y3zBRXSRviRxFcpQiE3VeJ1pANAnkIexR4xS9T3QoVVqHRz5Wj0FCMlk33shf2KJ
7JNRhyVtG8FZ4qi2FLqrkhVEgG937STvQ8rgjiqxXLg31noZziSy8FkDDcoHO9Fp
uABZhfhXq/TdjeYPegRzJMJjE89xEkT4pYciV+jXY/qL53F7utdWcmE6xC3s10Z+
8e+lQu2Ck7E/SEC+YRqYGNU7yguZ4JgKvuxi4LiPHcxwAVUAfK7sW+TCFwekOZAK
lhq/rgycikflOYhGdSpkloBZhOHce9KdHN43gv9Ty5pFFMaXd7b5uwoKQ6cR9aR9
1yVuaqqXXGUWwxfXIQvphU6VntHMpwjZqCF122DhV8ljLANKIyDMiW4kVnkFXoYY
+ADVXYZP4nwVE1YetVqJZb+d7QlLi5DmU/rBByFocXAPcZQIX+obIP5A4XNAejYx
2umY2uD66V4ZU9uD4bi2JVzQrp5rh2kbBdX6iz9JISfNaaEFrMY5W0s6ijpFUkxe
IDCg26m7Hm9qtfVsiKvNjWeclgjrWxSIJadh38Rt0NXNqi/E7N6ksj99v4GLWfFL
FMmsMlEF683w79HlXPO9vgJ0SlX2E3j8eNOxEETUsyQdWHYuzmVdBQQwLf1x3U4G
6zfTWnvachuwB5Vepmsrn97zPWZj8t0q2nRFXqJJg9Pm4pCuIAxV/VDJQOfE2kNV
sirYcNl+fNuGRYN3Wl7FKMYi4DZtB2xyrrqlCzA1PQPNG7fcd1T5SlZsb6izcTBY
fZSGxuZWexmyH2iS9Vdga+nqlZ0vm8TveIhUIhHFhqPXEURTDLaPMdSBavYHMX0+
LJdou6DtoEQt7YTwBT0iXMHkSk5FYrRtnBq006vAnF/1/96SsC4UdhrGk0ePHsZN
MpJUBXki3g50T4twgrmQSkWynleF+U1F5Pry2O2yxqdyn8mr/XSEP2RTbxEl4XQv
C2JbhQW3FNleLToK8agM8XppZm1tb8Q54lC4c8Z+FFdr981l9Oov/BTcr5GXqBof
m8RUIpcbTsvTc+l4N/Bt0k8E3E+Q+VaWypPYtf/FyLJ4RrJUyzAkDK6z+rCDppnW
PdfxkIAcNTfuJN8JDbU6t1seT71A3gk9FglgU+GnMpsATryBZ72C640eCB9oPxwQ
TtObWRDBS7oUoWsRYSmpGn5dULU1Ln/MGXp7I+aAV2ffBOXcZZQ61t1jDvU89HI6
D3LeFe70aBmsZ3wzn9TCYp7PHREHHPWnEJMHyYFfeWDSZBQw0L0Bq8Wnw5I2hvGR
mPKveunvFY08LB61laOksxz11IN+XuWQOi+1dSHuOI7eQ1iopxa0b8u/JvEH2Ch8
2/Gavqvh4jRlRZykdUxz4SmmCFdETy+e/e2/S1OJR63CSlTyQ58oxbVE+vz++Amk
Kbxlwm9ZlRUPZg2ca1V8NrQ+R6pgJfZJo9SRL6tNJEMuCqCKmbPQb0fmnYVPqr/B
Xe0ULF7nl20UlmrdPMLWcZGvVpgAkXpb5l5Y4eVvWxt5A1Ahn5P/XklrQKv396Tq
F9X4IbjN0xTsmQ39/72kYvK3kdm7XmkcWOfOT8m+UrMRIF3qe/QvAyaHds7SEJ/k
+bNEkPfkRcIPD1FEcn6oz4/dwP3MLtoERC2VoCIw4D4uaWPq+hTZnAolAY7+vy9y
uhNcieulWICT8zx4ItrNUK+kRCuzQb51TXlZgTPqmNvnpQD6rweXIk3BE6L5Jlj0
PNgnB5dfcJgFoX4MUXS5is8eD5z6BDZbUirvtOcbvREFhnWBaKzY2ESbNsy4pviL
UeLs4RmiJezD32CEr28aVwqjQaKUjZcrdsAO7/A+aOZYc9w4EmdtAAYqsDY3AxAD
aI7cZR3/3JKEzUtELcUZPqP+uNVi+wc814cI6YBGM6thXL+V/ImT3VgfH2nO7oQw
ssZKhYrd3MBtDOIJeWNTVW1jxfiu7MqRZwTTXjPDe7cwA0x6OyKAVftyGvIKyvh6
EY/M7b14xGTaXjdDoHrxf6mduLZybJx4xzUiPs/Un2gA9uIp/OK+6xb17klbVxeS
hqajmOD+xVgLt5OjxfHvX00HzzCQf5YpbsdlVeUqb17BGjNQgit1d343tVkV86Pc
jDvMWTg/NzEPcaU0us9/lYIoP2BBui7X2gu5j0cyS92uENN21GcdhRu6y+zPjE8m
mXi5RSYHkFOhhycZxr54OvnOTxC81rn+yuqH2B2x5sQB0188bZsZ2Xedz0eCTfUB
lcj+miy2qltB77/narG6NwqTqX1aQKWCjNXHsrGs5+yOOBkaQG6qo8SuUv2a+Ocq
OkeyX0AxBux5+GakEoafCzxmyO7Jroqltnpe/SDaTCf0cTOXZetg3AKdnfvUK8Hj
4/X3enFKhppnAfrFa0O1YBob4uyAQ7SuY9nhlbNndQO/yq8WWJLgS6da4NmbC9Ma
pGXVLXrAfmvJC+mQ1HlQ7NkH5IvTm15Jb5HXRBe3pHdqkvShRWwowchO1qDhiecG
Zo8hKH4+SyjyaLtYKQBZRVeLXovGW+vH8381CWSGSjLtXOxfdWoD1Sgm6phz18pe
991uSSMwifTEaD2y1e2ZWicZM21ppQUavqWvCXwY9eDUmmq21upNvaFqdb3BDF0N
1YD8Nb91xLet9CKYyLGxaVnUeZx9OQ1/kTj3v3h804ReisxUizna6T2rRyxTxP0w
6wp1ZXWeKPPspoUXYPjPmEXtQlvDMavAxXl/jOwH3uUCK8ZaLrV7w2RE9VGi48gx
8GsBzQl+xuI9lnOGlrZ+crHnSslNuATHcC9roL4mDqEO7F2CK1GZClut3HYuG9Ty
5twY+fBj2GQggCLqsC3WxF6DqvR/0PwuW7EfVQ8uCT92auKRhzk7AYJnpZFdLDgn
gEx6ziuqR4TEBm9xiAw8oFOWuJkSJH0gOdXWnqN6Yy0O9ZAQQjJq3L4XSD7BliAd
yp/EyoiKYCWjNfKbnMKjbeWV72LwHsiAoie8UamBcrUa/aNQv0nVB/y9GxLy/3zJ
qET5KS4hu9huISuA6Karj7PkyHQZcsJ17cFqhP57xgfkH1OHtZhupKqXYbuJ2mz7
7iPcyinRx1pLusfRPUMHOQ+wMZeyc4hIb+w4BZFW04PmsJWtmwb0siwJ67BrHTqt
3ggTvdrjlYSmXC3yaI7F5gpHN9c1hd3DvjmuDwuJJrexgPZZ3DJ27ZeYcpcohYfa
MrRMuDTnE9ZHXsmYA8ysgpDNbAKfd9gdKRIYLaCxM31KkSmyhJfwI05NjkXzDqJM
N+Q1AmXagHHIWQCtwdO8wZmIk50L1V8+IPq+KYqNeuKIAQ1zjPZniJNS00NEeY9m
znVmRqClOLxytQ9LvOtdtWB/Qb8W90jI1/tf0EzMrZU72h4xLSTdzVulqC4LPa3F
D8mkeHBNMjnwcw2yuWXyD1TYKZv9l4tWQUFkV5pNyX6NqDaUVdBlyviKBBHzNqBA
9d0YgIDTzR+qH6wJqcmL9r9Zg5S18r8NpiRZ7dBeyTbxFpetScV8D1mtG61S+IW2
2nXTsRfxgQdfX4dPdB8B7CSiVeiGoeDPd5y84dWmXcxpJoxg5XUeoWFS7ev/aRku
Wb8oKHs3HzGFyAWi+0Xo8n/cyKd0Ty+Cg6GvmZXYZ2Anz60va+1xpHgp/+9lJ1im
kmUrLVG9NJt/WByG/fENaYU3GdiVLStMkK7fzTEYea3L4lEkKFO8kjI8jIEpXznu
AMIddANMubJsE3J2ZOUxNFVTVo3DQdurI1rrWpr3aU4aY23RsUlx6qdXZW7nT0gW
DjVKtNbB294mtnIFjmiquTfKvVzHlIEMY26DrhGW1jjvY9+V2XnLghB6QySBL89J
2jrDtW8t0jYD+ZMDynymSkmqK9jlEJEUGuq6+c4TXppHcL3lwbJxr53nMlQE9f/t
FmcdBzgi5N5hrrNTSVjkqj9KH/annoIWz/apqn1IZl6pZzzrym+XkHf1Hr7pchH1
gq/ODwjLNtDqC+2K/wy1iEGcD7xuMvJI7mbRWU8HdNi4rwrFVrEDvhFsaJUI5eKZ
QaodDrf0iQQgaAM7o5pRURPyCTY0rJdzo+MSDzU3rn8wK2dBiPxNzn4U2ENTb5Ul
Pn9VT3DkKW0iDV81Wo8DL7aRwJOJcXoP+SIF4ET9bUByhH9VpXOtxe6r0Xr+WMo1
w/02QfsB9vjHyWo/yw9EUBFpCEiehk+FcIJuGHvjurU2cUkO0Bc01BFLNOpNWe7d
1rk2yG801iJB1NAMD/PeaNn5vPBNuUNfcHMqfXZUuKe01E5VwS0IjorXKiTe6wIC
qxAC3rRAST64dUAmz+RRB/LHWK0l3619G7/nTtZIWNXj+1Kp+B0QJp5F4cPG/s5d
vDbWFFXTPnW8vXlTf+bUd1QCT/jkqkNKFySKncvsTELbqyAY09CsHBuiWggIMl7C
JmIm+WNIdD9eW9o0MKv2mBFq1HZIp8OR3DNWh4oIkTw+1Am9Wx6rBeSoPwbtVXaZ
NyGppQ8kKt8miIx3fTmVYqqNzLq9VD/IijXJqoOiFnU3yx+r5wnGuDQIVzsOCz1+
wa5+WTfgnSMgom9DivntByFZ60xqGwLntTeJFu16w0rwdioQbfHjiVAHr55jaEmT
eXYGGJ72hz7EBsDRQHPfSWjkzLJ7CaHnN0bIFrNL7F1MhTvRiApDbDEzrEQ4X+gP
EeoHvVUiM6413XSdQckQmQ9KA6QaAjcrQ6I/P49c168FzUDoY4dQLcZmAg5vM0sA
ZMeZbmKTTSnpmahtjXD0Cklgotc452n66MHw5A7TsjKqT1UO9bNizdwS8S3Jw9Uu
P5kNOGjfh92NbXNHT8itbFYYvmIa03+lgNvXrzTZ9E5BF8R9e2D5dBgAdsI+88B4
Nm8qUqspwfQitFaFJiOyvpFpdDMeu6NPK84d3xD9wQDYYlrQfB1y5ys+8iWfkO1s
xTuQak9prtccyLIS/bAC/dMGX8LYXU1MUP+YrTClH8LB6Nycn60oyGJ37gd4mnag
XxZEGBHz5BpMZY/aDbh4zoaLi0KGWU+/yrgrrTBtewixzgbU3DfRDnDe7GYK3YQD
nlmgdht022lsi4joWQxVHrNxB8NeEX2r5QPvbh5C5EAKnlBnsthxO6RpydSZEO2B
gqRqzrJCE5yAseGJoXZI2nORHZINXT6tprU3cyv6SOOvvqcFNtR/WGqAaPNoiagF
pjteWoXgAeUibuZGt8u6KPkv2fAQY6Q8+/V1u2o1vH1mtDTpZiKqTeC46qgBIQRD
O5iN0SGAib+9vf78bU1dQFtwDAijnUjGOhjKsIIib/uBt9M5j/1wHKYJYnNKgMca
wVwPyzF4F0qQtBYsyFs8GXNlOwaj7sQAAknW6CHvBrU/RvZbcmotrxpto1ip7gRo
xcPtrn13/Rdb6SSg4f0MOtkQtfvrgNbHdvhHgWLIsnsvXRDrkoMPeT0lV2BcbAvT
S8o6ZyND4OWfGeEGxl+iAzazvcpINbaQYucM1gUF3X83Cixqq8w7F7owAiWWGjwG
WFtBvzcBcyqRTxLOPM02WHEVQhT5RaIEqjdwgLdloVLs2dUW+zzKuUny8ZPm75f6
2OisdlxeJIZGzO2VJhVPSCH8UnlSvUN8w0inLSWhQzO8zw93BitWXTHgk0WNJL46
Rvdd2u1e3/OmRhBC7gTg5konJED/LpsC9E7mlvOse8UWhMrYk8s5Bcw5lcKAswum
ZzeHgEKSep4+vwJE1PN4hWVYu3pmniQQPhpeqTFwOKNebL3P6ZDxIyI/22KuucZe
LZs26M3WHFqeutwEHFGv8LgAuxSozm6LZrRASUf8RmgvkOuRZ48kDLoCymJa0yjO
pjRgoBqmNv8ksw7AscRuv+k7gimX8KeTlPAHxQP6V4exKQLwFpH3DbD/sBfIKA61
GQzLhX1oeboCUrBaBhiwjx8l1j99P+a6Q5Nv9epHQhVvAhWpaTkRuEQIFO/MCsXZ
Q76W11R5mwHZqQn9arEYljfyDBXegq22Bb+n1ytBHnmgn8GHbJ+78NgOe+atQQ/5
3gXnzAzba1uBoeJzyDlaSHwy51h6ZMVLl89MUx7St7QDTntkdIaGwYqv8T3ZUj06
BrRXf548V0i6A9g8Au+hSOZZh39hllF07Ny+YcDjf4RyZi4sWoLodYebFfLMHAtu
A1HgPcjqF2Rq9YXwuC6W3VKfKhzJU76p3en9KaTgEFfo8mjLK7RvZif58Nk8mMd/
Z1VTgkveKsHc0ONRNLMHgF9FXbOorv92R9U37K2DkP7fqxLRtsCh0/NzPTKq3CY/
3l7WesuUISNUd+/xZiRcwhFE2+eoJAW1m8hz9Pyjmdec60hy/AYtyaVVAuJElHxb
tfJLupNZcGk6rop3yvGzyXIDHM1d5htTxnumloFd8LWWxZ4LRVrYCzqpyHG4f8/y
7/JWji/XCohPKQr87+O62k4ABPTIB2vmjcQvRgDVGClPxjkrHw5+bkhL8DOds+kD
lwcbwS9x0zctAegkGpffD/hMkCUmAYOSDtf/23/l374s0uOgbuWmN6bE9Ks7L+NK
SvP0m6Bp/nT3GfscrdLNg0LoHs5fb+XpyuHlhtgJa4j0fChU73J8iyBduZZoJkty
NH5Wwn3jMKN0ggB4CxRpjhpgTbW+YkkMOlTX1JJ2AkH5Oa/h6Q4OUSuLC8fyDz+I
YS7KNEVYTeiq50M8i8TewXoRSVMPVrFKH75O30qAgHs5IBiP0E5YgYGYyn6ci0O6
cKPgP+JfIvmciycrmhJ4HEO1GqjBB0gw3GpujWhjgEg3COFQw8NQWLdNkRQAZ4nO
o2xQ3u1ylBoSoxtVKvgv+uQZhOy35wCenJx/TvRBuYn9kFKGuc3KKXQ1hGXVvjmH
QgQ5jH6H4aHO6qVpUZ+E4lKebwqOUSwLtpTG7dPVEk25vISM4HGRRmyGZ+aHm/s0
G1dO6nSdr9rFoClSyg3QChMGVcEDiD0Cp3hO+eg9aqJh3EEax+Qi9LrHGvOYpUPi
JKmsROo9lFmK6WPEHi3efTIl3zfAn+F6Z6AItNOFDv083rXIOnMiHyGp9/n7/vCB
qvUlykfaJtTFz2tCraumss00ydAYjIOidIT4MpcLt+5/T9Vhye4mNr6Alt1gCuGy
KWTCNx2RVWoy1gkiMMwG62Z+qXvG7F+NZ393PV3CxVz6BYcuFBEAh4vJTbMzXzSv
83P+l/2IelTOhiloJFXvC3F4SVb4DZ7cZl5DPEShQp2AEMf1sDcdDet9VjsG2fJy
5TeNWot8V8gJoR8nIRoyf+ztR4w8CFw/mHqTl+PxfKlNq7udD8XGPvrMEfgJUYrr
QF0RwqvevlU3rmR/sOCZgZZFqIsBtRLNyXRc0KHw95VrppkBAriODKzNXeOGL9+/
gtt7088j8aBVukb7yB/vU6WBBGdmZzyEwGYpyX+ShfQ1VGXWcwWcAGMDiLKxAXcP
pAEGxLgZWt9cWx8qXdt6YxRdRN4O/WExTSS3gF7qLhrK0J2EYfZUNFVwN7X6DBT7
kaAsOrqW+oIgr8Gzi9lCKBQjWwhSVfjAmXqI2pdlx5VyHLPqzaLCpIoqgHS3MHlI
LFxI3t6ZU/uGt4QMDVS80Ef/4yw4dNAREsSEBj3Jpy+o/BqMCd7/rpRGXstI//cK
ryYFeODc7D4HIFYypEFTqWOiWL6jVd8cZbLfrL/2R8d7e/Vah6sfZasicXSlbFtC
0e0FX1+wiu1qSJ2qmzhm9dojmcG8RH5KvatgYD5qeVzE4SSppdW7L2xI+1rs780G
cEbpJU7AqGHh/tLV+NEvVkICOc/cOVi8R/0XRACz894bgdlzD3pHLYaBk3z9fOgO
TzgmOFazXQWOmKa+uPdsKtaXKEkzLomwnW91aWktrWAXXGUoegb9Hg/t/AHrEN98
Wyg8poDE4lqblr4V8CR5WwG6eddbYmg3KyGQqtS4IwaNCK9qP/5QxO7AnFmEsAN+
32f8VAeGWQEVB+rtlIpknze7g2PAKka29JS9pGATX8oLUu1Hwri2ZUeVwb2frap5
ZrXlkPcNTJ9D+let2vd+bUGJDrB6bYTLAYFPnpkjt2wOEXHpmwKZ6HWo+em8AtuU
KhT3gcv6svpqPzN/61F/+z1VmK9IRoREiIPZsfHuXeH3WipC4LSXCwHD96eiSrjj
AFCo2LS75xJdGFqAszD+OM152NKOvaMPO2YvcoUpyGOTwhTw8Bz4eMaC9zZ/UL1V
PNBB2shNKAbC5Iv5YfH0Gy4l2qLeLICNHxKIsq8ndFS6IEDF9m1qATR1XRFAL4pY
TJoYchsQIuBFoWuFCH7TQXrV6fRWGvf/5lTJXFtzNrihTVUVqsM7qzqdq/yMPS04
3i6QzxZIY0wCdRnpV8fLumzAv5X2O+6DdKbwBJkL2+yI8EcMWpiDmkND5BDJuT8C
PRkCzAqeFbFzw47l46bX9QpLYCzEH+CWAZYH/wJcS9vtazpbq85kgDk1Y2Cjq41O
fPKThGvhLSXUMZB6M+OWm5Qc6FzNhi3IxPJvkCvKc+ArZw1ENQ2155LaHDcYdO2O
HWMM69peEds6+xPZ0PATbYbrNY2cb3d+QFdOEsutKvTspVqCaQ6ggbF88GdFe5Cc
+GrSIpUfdF5szhorDVDv0ms9l0ImphMmYi8T/fO5oSYAhCTcZ1VJr23yPQAMfHiP
9FNuzm8igcmIPjNsJ0f/ynLRDZZBsyfZROVcIThAoZQspT+AiJ5TH6+AmzHNlyqR
+K2y59b3Sd9uGVAzIFgLxT2bljeunjiq8Zn3kGtvdyTGgbF+qb+17Ug+VXqWwNMF
mcioVuh9Wb2G/ykQgMCYxBcSOWo/VBDKpsRUSmVI1yR+E9vFQFwVeozGhwyzbPZt
4O6WDkrSvHBHrqIDcjYjT3C2PrpeM2sxioHiGVVMJFcIZBOIkJ/+KgD2lODKQBrk
Xax8r/Er6SzyGXkTmk84+AmLFih54BSEMfZVti8FEKrZSd6qf9LaH7STZCy1Y0QS
G5+bQ1vuY8+VU2KZeNOITHJswCqNZftSKEBXuJPhwjiVjQAWEnR/2JLsS9MGSQbf
wX/Fa5jD7bmLkGOCZ49LKMhsMwvBBC0I/Ynlp/tujV+K7VtSEENZB79hDebuX67V
BY+POWQnPP4WXir0/Zl2KwW57NcN8G05BZtHSKwXqeAcUZ41kMXwNNdW6fSj001I
4N4eAUi7DAj5ULLao87w7nMICdRcqYZHVLwvBuODF+7hXijdvQ1o4+N/c00z0xp+
WUcbFcigx4srJyihzT+9cZwUzIqQVz2DJQGPUM3IVrggFXfp0UENkndSV1aWJgzo
jO07fv+R3VBlDdn1RNAig/JydRdmG0IuRjkj6iY1FhFf3ltzC09txPynvOGBwAV2
KVFgPlSl4CtaV7L5nChZL9r2Ld0f1yA7537cHosKo7c3X8/NaAMiOWzYC9pvshS1
H3WxPE+s2nOrQ0Il/1jx4KX81wNcjnkeBM150sb/nNNELnQjBO26aehivdLK9sEJ
X2uBkQp39B91bLfz+HmjYcPjnOc/PZyloxbq9JZJU6g9LP7C4r4nvA/E25KqFbG1
tr5cf5GQxTKdVFeCw9M+Kr6xn9UfZnSzcF8AHtox4O6mDKSWK/caHKKlgREQWo84
PMOKRJIPpVzoS6IVCbWZl58q3M+D6G1oDSBuw8DWb5dtHmZJZ7hODsQqIUaKwYQu
vmkwwJo1nXtGfuyhhnTLYaBvmIdSHF664dtRu6UtDu9n8ojITpODZKegc0k+1mee
aoq09NoZ1Rp0yInvQyxtcr5HLfTitcYGIjyXyeiN1t5sGBv6DAS51yzCQFGA8jGs
NkA1l9tubcpp66BOZypBpHHJQPx2dL+st44F78/lbmRXbkAGk6PxYzXD3+rHce6q
jQ1W854plJmCUIp3EGuT9z79B89Ry0DJYgVrNW5L5UFJkQ2Y5UuO6Hfy/zEoLS5i
3/rl02pZOedmAItKnBqugoZSu9s7Msv3Sz9b9p0jXbjiEAVtcW8V53NCfNLZThqC
xpJQTeoDvsYyLJ/tSHa/BQ27GhqxVoYID2DIksoNWGdWKA0LbWtjeBH5iCcOb2er
XhxGHmke5DB/Cf+peAcSMbiHgiYAdDWAoNL66U1DTkbmmPPsvdV7FdoWGk4i+vaK
Og1KiEIWnxupFfh50Nq0ldEUikqiW26kyHnFYSUbwFdUiYsrEVbfDfhw47MpBqDu
JxplDa+CHTN/FLniVOtLIlTMQX8BRec+0ubu+oc0UW8sUN3VuJtqaSxISvnp71oB
RPMabWKsOG0H5AE9u/kRtw3ElGobKfQTcH/XzfiEyF5SSmMrHQSZTjYuU0r4fwRQ
2zO+zxCsGhRvyRx+uICfgol/ETmI5amNlSAN/qeoIlVDqsO7C4Mxv799bzlrm7Qy
LKu3ZZoGOOXzugZDs4Yrr+8FnznfsaerozH8KIR9O+4FV2j1Dcm7xCIgFo4ZPEKV
OXBgrrExu3ppwadEuFnOWVE/nUtsbrhDySem1oocahosyEnutd+ny2FHjPpW2gUJ
+tu3orC8N//vHkU5hbTgXmNtMeo3gGCD2sC85rOtqpilSR04T1aqNJsgphUdlSG3
CifNYVXHwYrA3DMY9D7rAlpGXuO/DruqM7fyNIbHt9eYLOTqvfyZI5MnGM0J5kU1
X7wF8rvnfpgW32cavNW/zyuqwjw1o4zzpb/7bHrN+gnk1GtosX6KHxy3XJKqJkD3
RH8mm8ixuNngO3o/dDoA5aXAhK3/Pq5STr638a+1cqKfEh5KPrBxApAqJB+jpbwu
pUGsyptLuJQjQzlN/ksGvIeie6gcgaKUl+UeROom/PorjWpVjep6EwfQMxwJColg
KjI0PR6QdCJfy2Om7uR6L78/KTB+G5DzEcabT2AzBlH2vdaMoxUd1YS2oIvFMyGD
VlENlWIuOBQwkZgN2JjRffY0ycGM29HDBFYs3uKsXooZ0Sf5k7WwEXotYOKSfF1O
I/2G3I19lwSphxe9cYkNPrRu7KxxT3e1+DZnB2kAlZRlxUUYgiZ4iRqhePTSu72l
Dq7+t8qW5DcElj2jb5iFLV4HHs8nGwdfsJnjvEZS9uAelgqE07j/b4Lky8vPN+xm
bisMxiLrgktMJyl3mIS5rWLyiUq+yMReJYza+2QnA2/U6Cze0DIeGj3AjX7H591V
v3XuYIWRBlff/b4C1Be1KPZUXN4SBT849GJlP3U5YHVRZvE0S5T5Itqvq9cbMjoG
v0L3V836+wCqYl/VJ+E9kFNqwaoqm+XV6p+81J0mMY9iLTyJuxK5TLGGBLSUECT4
N0qjfQ1DZHuFe66/F6e3OC7NJgmBMamJSce7ASHh/uz1aq/sQMzevVAg9/WmrcaN
SDagrFjVJwDAOXSQZ+NiLjVzZJnO6bv8BoAm4OsV/dEOM9YCOG1WJD9dOpC/qYZA
zOjOtSTOz5j7v2QKnrQwlsYRBmzeR96wEV8nLCGz1/E1r4O6jyG0JKMfNLFEOYCl
cB1sIpmJLuWGxXYkKpY4R8yAciArv8OrEoDW7SUAdwAu7LswQP8lGcqb3DWfOitp
7r3w31kcfg8f94h5bdUySxcjpMN4QiVxBa7RDBGnQLSl4TG3rOYy0HrxHQo1YIIs
fPGsuQAd18OkV6SggSBhiEEP9CVVmwZhKXJkhyAkG4JVdMmW+Lv+q10QPd5tcSDf
NcddJdPPydFO7/VqrkfjCRYSA/a6Gs+QEZZs6fZJmUO1y9v6VcmSrFdMqsk09zKH
5LvjuBXfM/KrkNiEwlLYARqnNv4Cw1/MR24rYpK4/ymaEgB6JUFlh4rQdYhiam+9
KOmqrdrWCJ1rMYj2kFnjXzyRv1HEeThhnnZfoe7cNV5UpT5EsADPL5bhU62DXpsj
mdyu1J+XrBCVdeQULKebGM1ntrJCs6smPMi03NLY7O1OVt3DeC8LHSzd0dBMCLC3
KAXjz1P8juRmD/42d2FsBviYN27hcqrQgEP1FM87CbkrCRWewqlVaNAQdmXoKjUw
r6UqSY/E2LSIVTQGdRpz/e0d19KoZFHQA+/pRGXDFndwmu1AtLMscMoNq9ZH4Q/W
CBsFFSJqReRv7ezAbMj00a9bHFyEsbDxlpysADTzLG8VoKh/Xm7zsF+d9iHYTxLI
CkgocgCURvqkX84T/DEWAKKsmNRAWaq2r/mmTzKjue9hT9qPhisOZe9QFxRpaQgX
Zw69MC9MGP9CU078Ix2N99kz+MBiH0xRAYIGAiWtyvUY+WV2po0GFNuUAGWrCYoZ
ROD1EkG384e1pGKtFCxdcdQ1EdB4iVNT57/IZK8wF44Lrx/8O1dVlHkTFTtq+dRb
oNCobfHJHkNI0wClxqoPzv/IRmNLxWaKUjirs0GiVPab3AewJHeHWBNyk+1JC2Un
/s94Q9vFHZYAOJLCgm0Q5QOAXpZ002yQhiVjG+xdhZzh5jgBlB1ai4EtRtRjht19
ROn+d/7y7Pl0trVWOlYsMgfA6vvbbvZSo0+r0i0TGwJ47Uwl49oSjTf3HlEhwyeJ
76eoleGdfWsxLtxxHTmvQNlV17nsZkSwv5BKnutrEs2Aj5iIZKQPEuYkCMJrlB5a
rdV+Sux3ZROBsQXf7SxakZzIqLjHKglbWP7t2Sxn2lt4rwc6Go3TaGKDxXm9/oaJ
zClufiVt1BPn74o+TSyydl1eB9P5rQwWKExdm1L46G2qrDhXaTmX6hQI3Ofis/vu
Z04a9g0t0Cq3fy53tHc/8146vBD995uinuTG7necLSW5Vqf9Ng1iZrekzDFatyyR
8zkiDlDVpyk4sYYRgVQChRRale6/c8CYN7u5+rDprgtMTDr5QcnpByIeIA4H65qg
izROP9+/48GemiO7mRDnmUDrm5GRuKaAlqaIJlVohxaBgWOV20BgtNt1K0UZJMb2
qYeH7j86jZYwKGtp6S9FoVykgVcGu7BLtG+FByfyJoqY+T+KpMAb5qQPsJmzqF/W
ya4vxApMEuaEWy74Xx44S4RBkz996dovWqc1pgejUU3dcFzjT5qs7Jx1U4qfJJWu
QSnaqVC5HuKq19iksqBwBH0vUiQyU6NGgB3331M1VqGntYrreL3KkgWFMqQGbTaE
GIS0L32/gBln20a7wOyLDF8AX2a3UWhShaCTCce8qIaP0z9PfeFqVK/RJFcZt7zM
ah3ApwLcv8r81VnfKL4bYvI2GiJn+Hvv9CiuEG1NGLMfMDV/DLFz8aqQ9ICNPIod
PbCIAXcJyTxgAZE1pqyqZGnL1q4b6FHljWOn+6NFtZvpFGBbwF3SGdDMlxG9RJH+
uZ0FurVq6V8EhHWqZezclQ72WPb/4P0MjPOn0ctb2m/pzR2xdZUl/a7IAqgfogoI
MY+sL5vgnW2yU6iIQBdEltkDWJcVn14/lTZU0Xw3i25vbOJDYiY7aKTmk05YXzSh
26cPMsANs8xR6R0C2GfZ5Z1kIS9jnKejDWhhdHonPnxGMv52oxFuEnenLy5enn9U
Js/VyL5Ac7ifrUebg5Xhxg3/H6BaFTlVtOCbDo0QTOl6YO5+1L9OJhAPmg1LcdWt
iPfAB2U0j2wROFa8A2wT7DV0iM9tNCg1AU6z6v/Rv23SlU+gi6TVmBqrTBO2/FbE
yhk/bDJQKfpwsNrBXipAauhd9TYC5TynqAeZycQZNvfLmFJd1oyDX83BJQVAABko
eBEPzzFy1vS/zpm+qlxlEq2s3LFEg0V4Af/kAIfYKXFjTGMQ+I7TdcwgbMHDlNL5
Ejj7THujVig/JPMU48gcmXEQAgOsydpSPhy/M8x7ogzmZxx/n2T2vzz/bnqHAvPC
85eBx+kBYcMHal61OGTadsOwMexnHPE8RQUYzAbcqNVRYnZckmksnZ6zTYF/ck0Q
YSK+lSXsygNQFklsjGzWqzYLFWwYSV1Z8kZeIQJWoNluuVXcHNM+yXz3RDjy4JLo
bJ5GyuaBWR9Xmlv0LPUqbl/e3QVZDnFJSiKfbX4UN8LC6eDlr9gX1pG1m8RxQhYV
cZFEHxpDcC+j+Ap0BUsazTPwflqW+84/g30aRjHorpU7GpIhc8aGp4XymZtUwx6x
rdxWfhKbZXMf3bBWOBec2KXhwMPCCe1tZYV8+nIXoZ3K5LvgUFUBl3QWZ4KnTkb7
YJ68m8s7EeOken1hB7E5PA6mvoKEteRwWyzzIhIbefom+f03mnXYRn8qmtLmBXff
fs1vIy1ah2FCXinJr7l/6lHR/m8xPTjJxZthgg954DyhPl40jD8vEYWI4h06iJPW
VuSkPxgiDaluvUtxUI4fRtmc0VOyU+iqv4SXg0xDxTA9P3VPvWKMbc57AGYonz5I
UOUBwZL77CRu1PwYyLBJudr89/SPTZkt5aeIxFo44fgN+4pQqUc0K5o91nTNoTLF
NHikSEmbW0e3C9I8MFTklQNWQWnPpENgGjo+m9oaQOMztaBmTIGp1tuTBnJF92R6
22avkYsBTwjjDwNCgHbV5zrjWM/6GmM542wuWOSPuFbBbjUMYZt/SCq16zu2uiTd
VedT1b5WzZQrxOv1Lw5h0pVJpMQ8GjKfxoytrLqdAqtxkeLwK6JJXso9OM4isQID
S5kVTTHIZVJh6YHqeluNNXq6kjQQmHhjDrnwwzJy7k8fTpbQ6S9jh3GfLG+qn4Cb
LZu7BomrikaBorVYabia26cU8K8N7VASizWmRmeZC2QKstuIa4MTvkLW0ZSC43BC
+B+FtgkHveegVKLR/wiwxYUzJgLhYES15QNgmztN0ipwzcYxK3nDYi3RgpJc6jt3
JGv1j8E91EKxqaWPIHRp738+nJOr9583o2mv9EDrQbTfsti2mcbtXXuERAnzR8+h
nkO0yhno6FGSTWUHVJ+9j60vCyo1yJ8WWUY738I7y9LfiMYIF+7ET35KfokjLDuM
Rs7HW6QgyihkeWHojx+uwI1jw8kS7ZoJiQJO+8x/uHddClbVytON6gV/M+n5eq4X
85wG4A6qSxV+57ihzxTnsuayEba+1b4RjVwirAH47Ec2ziswWI60kMoNz5GVvzDp
+9TI5ArXaGqUPYVQ+txxXLMHvDcebQ59PhQrF4emfWAe81XgHE/32UDzeknV9n+Z
wtUQkymGbnTCrRKz6g1P4VGngXDw10P9zRyapEsRokewA3qkvXFByAkQHDqsqHap
K1s9+Ob87x9KaFrqCjR8UV5Ly/LAKeL5IxCdFDvx3yblbZ7OZQOypBTX8SlVn8ld
krKPka79YzjT/2x5HcPKVPd6ynYheZGeIyXLSFjvibh/aWKyP13cACWwJGGcwX4j
o+gvK+ZPyEojmKki0os/Ov9myjenc5VBVA1NJzNqTo4zHVvMNQ5vXPppzBQpSINw
o0gZ1S5IAyrfHGvIb57phq5r+bsBem4stI6sAuVQAw2dmzYAK0xVrwIryQiZnFOB
77ymaiZD4PhQksVSqsZ8xSQ5+inCSgZIi57yTvtofUzWAYojilQA9Wthz8q9qtyy
J7WjAdEG8JBKQrrD9oqlwTBGgylafAeWycoBDvIVnTQ36xBcB0kami2WzUaEXWsi
TAyRpzfBeDtftaxUj2hVv9N/IVn8jsxV6xWNBp/xSqcoLEF6FDscOuDcLGox4m98
9nrZRb8qDoyfiLCYiKqov3plVxVjDljZngj+LroLIar8dV4ti8UPfAIW2cq9amsj
XA7jUMVk6O+MRZIANZJuH4T9pexOfJurrLJgigUhjWnVnR6ReMKEirhVtNXWGQRR
fsqDEilncMzygzr9HdmLtCfqM0KynWCb2usphzuDMbVn3REotITdcSVlogHqBcVx
Z0Y7GeVaxjlyyNUgDCWZKpRNwZqPOENvQKAGowaJ/2621xjyTcz0rWm0PttBczES
Q57njy2TDx6C2pvSRU2M3wxIXAJGtflkVdQPWkjiBv38S5YbtFuTomJzz2b17q1W
L86btnKKa45RvKLkBO01GRbuCV+9M8LMkuhXb1iPT8ZbHiKrU1+2JVmBDVEE6/I7
mEmfmvSM/i/a1a4C5kr+Ut+01D1uojhFbVXfjL98qjZqJxWDfvdMwiY1kjQrGfSu
/x6Z7bkGNwhXrBQKEJ3DNZ75MdGK8XR35ubQiqjbnYlz9Q604znM2+aPxWgS++tG
lW10c1V/5VFjqxB9ZUSMeEUl+WjetGKa85gPlEw1OrpuwXd7kfL0TRMBBEnoSlsA
JVsUqKzdx084XdVEbUunOzaWuNa1eRNRYpvQMPvmcdJPEA1srvSY3A8i7dCh1Mxr
XOungaLavhMmSHtSsZM/G0axZCLPoRHTSsie2RM1xXba9q9RR1vBdmaK2BTbOSbe
SQl1edpbRHgV0AwBKU81+lIvjO65PUxOmh2WEbyWBKl4h6CKZoYh4BEnzoBrww4Q
4cxWn+aFmS0uGed3te9NHeeSjTAObMxKvVpXujMNbaRVpa8ea+q3ohxrhhv06Ctj
gfqMpBzzzr1E5RiHKTLSIlO2LownCSw6W/HiHeDpC9te9pOYN2FYE++izeGYam8E
LKKbYJQXUioiKrhArdNnDudbjKpXb3ukyx+d4V2Dh2lBEJewgNy1jBkJWrl/yojd
WnUlvzqhHa8Nbp+SD2BSdSNFP9Y6Nav6uaLG/Kx27IWLmPp5c32SMEGUeGnVPjPn
aNxaNSfOgWHBiv3FuG+zYndtehxRFk6kZxPhhBPaH9I2aowT5q1VtszfTO3ZM3kh
zHlvGZE11X7T3IgExjsZoTVEgnP6iKdYHTy03DX6HhWQwZcr5X1vymKtzbkd/K3r
+gJ87/H0ANbNP8l1VvxC1xjog7dwlv5iN/HwDU4HitjOHeo8wF8cYPqFTSVxTSbF
JLVnf535RbBnV8h6GQFQguKp6gI4syA1zAnwJT06FfBUtzILid1J6vSGXjimROe6
juvze0EDEEhlptUFsbuRJ6uj0ZO7AOZ3uWqqycRTr4pu3uBRfOUZev3Rn7W60x39
HD9nbuMZFH0BJObwqfgsiF42GFOENr7H9Aid4H7ilP6QrInqviftknnigm2yntDg
zIqv+6pLEagybGPLMs1naev2e+MFlrxOw7iKtlqu/2hHiuzl3GdnGtg+ubql0Bxm
OJGXtn0IW6HIKuDYKPL09aGyRrXgCltfO8AItQCj0cMWhqoX9tQSG/p5eCBcNHR+
8RH/koG9rT3j1OEFScE+7Bchf2J46G/zX3SAEfvfw3B9kteoJN8hHeHS+oXbwlEh
Ja6b8MfnlFR4seSVBYk3j+X0Tv8FS6Vz/IS8t5R3W1f4F0fK5xJy/1HLIz4Q+VX+
pBpdaETAJiFdyyHUIZNANbDjloOHuL9T++yYqt8zY1dQAxpctL8AMcNEohd5d1ZU
XWwYBi7OAXB4EyP4WdkHCKGG5hiS4TglxfmRuDm3+2EjzFK5ndyc3wDcnNoSrrRk
dD+9rk5uEiz8kyZEffCn8JR8+YN2Pe+2HMYBTyFLBq+5rP8fF0eB0GdlD4tgs+GW
yVVf7GN/VNBuVJLHGHhaJQo26KTNNk1CCh0JV3fQUyZQxHGUz+0kkXbEVbXZLKBJ
83dH5+1FQXyYb9KOajxpdfhuTUT7n15H7gKXtDENAdfgmHnsOnAgNRCdyBzkVu+m
xtb9AI9YFoOjKPwLH9WbBMvsgMIj6zvl1dnMd7wNYk8AIMRbyBuV8/5N8ZbAGv1R
+tPt2Pb8mBXjSCyIrvG4n5LaFi5JJXp5jLwGytalA2nVyXKz1ixxEWkxJlVPVhgY
abEf9E5DOAATj561m0dW8vOtlZ+/QCboHWm1w3Vr6zmoSpEgxjAhhoMD3uTnLGAg
nd9iVsnY5uPwaUu1oo3pjXl0BojuBJveEIZbxonTJ7OJokgGAQu9Y7EzzfzWMF9m
mnojc1pmoBUhJokQ8nHgR7KcKNX7OjYtPGmqhFxCNmuOxyFnB3VPU75pqS1PJ/gQ
GOVQZk4JluKoWUGM2/zDeDz+4y50GDCINZE1pROpsDA6ZV897N+x2FFo3/j8FaSL
HD/xRr6YKjDHY12/nY/BokKU1jEcCSNM9wxLewpZKHRZ27rrIMX/ZHahkXCR1DyH
RhbNshvcrGiFYZeQXJs1Vx+WZ4bRmWTiWWAoshmF50PNUUpOVyCxElxAC74Y4vyz
ZXaeCB94SRV7RU0ubglC6QL/SHx/ddq/V/HRDEQ9GsExiCWM2mcQ9jutlv/ghL2h
LPkHSFOPZrAVG0+WTGQdW1nOhneLLkBH2/MKs+hp5m9PXJQw47ALzArm4tjN/j4D
yo3Sqh9Varu38YEfgyUZ657C1ceNlY97vfyAZUllfsJ6eSI7WH+BMGPpJB0c9f3n
zI3Fq3vGks5g5u6hDVj8xGwdHUFUFMkEwEOL9hHoxBAnzQCKZFBzdXD+Nv2moJL/
JL3pBMwqWPd+Y1UqWrLTVlelCf3d0y+GQ7KqY5YlLiuWboLjfH7cmxolcvJqtqSi
bShKUgp/j6pzXo8M07yQf4leQspf49MVqQR3b11QgEDtiJ9r+igk11bvxdmznYtj
NmDrSq6m7hOI6BWoZymH4HIAbPfWCDgtbB7uAQQ57OoydF7SA2IpxgltBSir4SWp
aBeB4Gi5Ki/8HHY/w8HnpayWdwEEHXFrR3urjwHWgPKacH59s/wVNK7MYNIZuQDV
TIhOECNkhA3e7zUUCw3/eSBJqgSC3uOI5q47z8W1mIC7FyO4OPB7oNvdElVrBQ3b
yxB8Fi5joCBQQQddkmBJM+a2lqNwrUvL0Et2dzHogVPXggcn3WpW8NI9gwUrPL6X
am8sLrVqQMzXqvNXWE9x/k5PKTiZrPhuWaw+LTSvB7SPQrJNgNMMOP3QDHFgt8Lu
EhHKs8AdP5qf/fX7nGuGJzPXYhWSZPyEVdkb9q8lvJ6eSPZ2XFEBKvOkdvelPmFE
BTAL7KJXnUMu5ApXw9mETlqixhA9PapcwM46heBg+b7ydYQZWhwv4l8VEm+CY04W
4Firtg2Yn9fWBwhPbQkzWqK/ANt37i8Qmqrt3OJa7gzZrr1XltSHpMqf6XeUHsRn
dZlpFTEWAvpXbc3jb5Ruk/T8EMlYy7dn8Y5ifs6RfOXbMxOb3MfHamYq47dTvXFF
79XXcsIzOHei5LXBcaIbUAk3ebXr3qAIVMmI33jDNR7pa0wgQeYu0qx0nyBkdgjM
oH8ep+2t6SNo9aJIk4Be8hyvJy8X3kucnBd98/EZL6qSYLVq6mevfI0oFli17Yse
pEW6eQXitZQo5VfRVsiPEqw6dFfgbQqNvsINB2mHh65lD3vxmB4Mdpr0Ttbu9qAa
C5Ujrp7hK85X9xbQn9L8u1q8EhXevmsG2LZxLmE0gmWtF6zk5gaL5LfXFmq1KwqC
dlJl5Xjp/HagRtoFaArlcs52yQ6cZzIfX+f2uenK7Su1IOSXzrei6D719h+51kmR
pCLflysnFXmGACgzrNaQRX8aycRk/Afv1OqoD2hMPE3lTtu6FOfD6ozSu9k+10V2
GtSKjOI7JI/JtA/ma/ucMyhPtUIdnBlLRtGIkaN4znNvsp6q/9YsN38vD2L/RW9D
TUaByXKehmTF1KUO72gFo/53drMCsCd1u7QvuN/iHAg/JMya9wpJYtChYOY2SdV6
n618rhkoiolzepb2RRiqcN/9vyTxSI0cS2J6Fi5RidJ8slzixDWUbO1VdyCG8yFu
h2FZDy5NhMpjkI4mBl4W7j7hyiFgGqLMNOlmKo1bjWHiEA5xElkLs/2xSLxz2nbh
U1RrxQtdhcGjdYhIuL+RE0MioEVysGbRrNa/EEFhcIIDqhDda0K2NVd1T7vNk4XQ
gQpT3jA+l/f3IJXRYxdihzMRs4eWl5BjVF3Ew8+5k1Glm3bGBPNGHgQjoS4SmAuL
ZDgcAloHsd2XnrVuvPvEYbXPx5yeZXFJmWZcuQzraupIu0btLI3XBdPevf39Wld4
pLdhqAbVqrxP8IM3q3XCkvzgxCxq+48zjfcXpvx6DGuZKZovMV8yCZZicDiFXL21
rbniPbUl2ccRJlsQBR02sHLylwjjM5x/K5a3CHRkPKj/r30rccCHM44n2HVPc1c/
9Rn6cdLZ+uEq7C74EhkDpEdXzGPwF5Sn9H6ugCMXkChSum/YEyCckB0drpmTgiMK
6spC6Oc6oGuKhrGdFFPOa2CXxAoslMsc7w3tOKq6odQWNt94iZnuMce+VviTSRir
P/pT2jrRM2spi5487vQ6s+hx9PEaqvbJtXUkoUO+p2f45XlS8k6pJm+RAzzXq0x4
VzJhOicwChR++tQdpQ6hgLYoLHEW1i6MSIAsHQi6cm9xHIcRxzUFelqWnv4G9aLo
KVINtPf9PsoDfalEHl9dLhdyuy/LLbwhNHLxLXO4uB35Tl3b5nS3epyRxttV8/99
eomgmMIyGvgYO3b2DIOLp+OvLuVjZNzdi8BZC8uDu6G5sryx5AUVy+neq4Te2W08
nPQ94updttDbwOgUz3629yaSAfqsoacOXKLqtMd8MxBsB89BAhIsPBb5IRD2tlWq
8fawSQymK3f9MUemBNRyg9oPlNTmhDyWZV5BA5bRjQGPXzFWB3C/hVNoBuMe/IA6
Ak26uROqiCQ8ozecvxFrX+H7WpYRYyYusLLeegl+wfHGIchbZJ/AhJuojdPFz+US
4rR1XsPkzglChFIFGB/rqSA1wlUydn2DjrfF+npBgKIIutoFsGxZrxTzkIUoRN9E
2L3UoCn399ipLROep4LD7+1r2ueNkSTISDT7jvWgFLnvnz7/m0n/OOqresS4LRSq
lxQQ8JXup29XJchPIGYkdhQzpC0uHmo6pnhhX3Tbc2And9hYxSwKS2M2e+jDJkQ1
P6pLLe8ZqoTGc0Eb8fSEcN/r7EeRoWLLnGmLovxrR7oKVcEAw3Tzi7OPVFDYtVl3
HN0AUWtMqUeu/cqiPzbHcSOWyCyqRtbekyprIr4pF3F+1HUXWblHv6EE8an/aZG9
wsY/QSHp8sB58WPiennpogeGmwhFH5BfSDI4L6p2xVs0xBd55vyvEkiNs0xIdW5D
Z8ZnehMflF1RReyyH7/XpjjZyV5BIxDI1XaUARLATZ13+kDG2wplapVH2nIDStuD
rjMBeWLPGsFkmqdXJsAChuX669xD8QCzhtmdR41P51BodU/Y2JJ/EZIeHCXjBQBW
kdsePyuubhWCZ69lkuORaY5reVDJHCD6BsGgOjtnSkVuNyllRBougpJ8HIpJRr22
qv7ZhYsCW7i2JSoiRdGbih0GZnHW/KP99Dks8MbVidCumj4vbRqDxEErQgp2R6wv
8sNa1XM0Dxw1TJa2k9Qz19wlCizReWCaRa8UJ4O5qd+c2uIcyWZaJSvIC28zv2Nk
M2OKGsDGaI8p7asx7XSKPx/FMMrL1j02RkcXUz9c4CtwA2oz+mwSoZOanppxjt3R
YQFjhEiZ+i9jaDdgZVTheGJtUZQI7Nn24V8G8PGD89ymThCm8H2sW9nwrIqzueoU
5FmfTV9sjm15dIBfMqqUKqrI885EkEpTZ35N07HauntOxwuqPlZtSvIVhqqGDtpR
GMP87Cmz/kSvrJbYIHxDJNAQlH4pd7b05U+St8aTicDCHGH3ndB0I0q7lH873lEl
lX6PdNcVGDhd+DpG8VklsToXqbUU7tnypgTot0BWHCPgP4ScVRAIDO7uXrLKEO1l
QJ0izVOc14E0ypKBcYamHFM07QkC/WLq+kYvE6WKrW9/eGKwjLqUrMzwlgmbZR97
e06eSlYB58H/Wh6nNOFrfdkSG/tgyBfKN+AAf4evEbHa3fQnEd8ZmHGOoTsLtd3I
CbvqzW+IMtDcHQ1py3cOK83Q1Gp0bYDGV9AenWaIwAPGQzUHjlTOG94AqkTSizwT
NXNitlH5KYpDgU44tDeb1cwmgoykz7rQIg5RVvsjJi+I+0yOhFDel+g0cIBxnIzA
LVu54yhi7gZjcocSfV4QsDwWDXtkAIMIiv8NUGJD1fSx5y8X6GEF1nyUi4TJzoLY
Ypa5Bin56fKPgIW9OvkmZ9cXUG190fzSmgIwoLLtP/lIxyw5+hPfirTiQO0asZes
Y7g0dbm3MB5xsFlmhSzFVj9cgzOvrulXo6Ybr1a8DsGHmzPW3tPmY21L82YomyTM
yFV9KJHaBZMSELg5SgULGQOp8+lVpbaNO11oDr8qWKqA3rAGcwljI1r3ew9y0qR9
7GxNA01SkTVkwi8mUu7JI1Vt9zvKLnfaYrUKhkPAL2nMOyyfOUb6JCPUkYnUa1LR
bD9abO1Qa2X6FIPW3HriTmUSMox95QsfWpaHWHTsEAOyWehaZLCtUNFeYkFwRTtO
20VLh5W0GLUOJgoAneZjhHDFEpLK5efebpgG7aOyG78aa9wDXtA+NmFKd9KfCh1w
XDcTfD94KsUPLjP/JOnIGB1RglKHqvjyHOOk3Q2KrfgF+r9bDJDa9QvA/YIynJVo
YYxklL8Q4/4RCIwMSxWa1+YJXqu6cOE2ncHO9Cqby1TMbl+YeMbM68Vxzch8XqoV
wsUe/L0czpntv4NDlGMwtXWICSzHn5/dSjnCp1AvMNw+F14oxHym1VSGYZVzAOyw
J9y+A234WjcxYtAQAzIK30a99k7ZcrvuquDu9+u7sKO827/wfYaQM8vw9TPjT77+
HCSfMLvzoh/wnNxP8153gQs/3OkRKs5fU++CnqO919K4PdbqRsiThFxDrjj9pgxC
N96/L4dc/EeUYKJyW1XzrH/Nm7hXzns5C8r3eFhuVkEaxWbRzeCYtTTJsL35V4NR
y2JUYJDBG01liMlIBa0iP3HRzv7S/C99RQncuHQjZRjxM3zso2KJRS8RHAkTyUnL
DpX2M0CNRj8gCt8BCp5841EB0/ow3GOfGeQXKvq9W9v894pyjPnN7XcDMX5Jxz6j
2f9TKKvroqzI9KgJvo2nKdWW5XKmql0lVrWRy9NePTKZ4js312f83yQakNYq/gxw
VrJoo4+sTzgdKeZ9KlBD2QSfeUqWBV09SuhGtBdyOapz1r/UsV2KvDaua5SPuaDu
hP96ZCUTWEHVGPMs2Bxom+epzk2md17NiLV7DEeZAenzSpWM4no4v1eqxZYeoDq2
t6E34CNoOo+5UYHDlDJ3qfCGmHy5ss8Kntwi/2KFXSQWlOop5j3bF2GnjkLaKjbp
saUNEg2Y2I/8uyU6zpEKj63KNAESvhLUbxkoBOCqevc3ct2INYeQzz5F76Job28A
kXAMZtF8JRsJdJY6lfCr8T/evUjFEgTr/JHdBypLzSBXo8Xl/OM0hD0lu57Abw/j
tVyIX5MPHQYGBucBJk9Ls1evSQck+p0fm+nLerVh4DCJKNA9iGRvmqTgSP5OrUe5
HE3VKpk7NuRRyCKZ/BmY86rUuJqR5YE0WSruUzcDMgkcTRCAo1Gzi+9+jijJThzh
EYm6G23NpMeBSYokMPp5geuOVrpodSTi2UoNSO6MNEGFjXU6FAAiHJYReyZ31x3A
UEznu3ZiPtXAYjF9Y5RgWh9Hls8JWpk4+VfrPJGRMIqAAPc9I4HhD5RBMq191mYw
G2aDntnygW44MWEY5tY7uBlbQTDMEX2sdWwmn/aGC4dpEswGLoBIOx0ltBUAYOiw
F0hGoSMnIz9hwKCETZ+K9OoswzmXxsShK59TDfaiTylWq9QI/U5bt1HgVKrfVb8A
18UJzpX87rSgKTHIe3T6ivtMOHG6A5EMcBe4mBumvbut+LXatk1OCu1b3b0VuMs+
Ofc63eMDhDpo8XhBbi/uIoKcCxaJ6jqfK98Rkij3HbLVexyhOau/FGoCV2EhRdCi
kFE9yq8ZU/ZyzRGvdOyzXL8FichRXOVTh/Nk6B9HO4V9LM4Y5u2U2tdqYkMSLTkV
ummtq3r9W29wDiRTGdGE7s4DFeOx6RAXi5pAg9jsX0990g/x0TiDa+PFtxmoiL8k
E97BDGz0q3x9WVWerivqfeYiOs2XhvVHE4itZeqDileCV+zoVbkuGeLdvrMFZ1NJ
Y5l4H+IqET+zIMXyNRDg74iikIhqVyxTOf8FUBeDessbYj1gif9pDlHdlk6ZgVon
ZndMZ1kypFGQiJM0pzJWKQ786m6ap40mnKjJNdZpmz6weZfizBC/MpSjQLTK7+WN
v0gkWqurGb1H56LcLZ8Dy4S7K5taUWHjbhH1QSUQ9Yh9D4Eo31DVJ6wBFnjzb0ww
yrl+YaJK+r4y0iVek1mVv920snIEbxIoMQjZgCebE+CsubEvxx5XURljvWYpXHCd
ayieVydRJvPIxwLiY+fpT2La73Fo9Djo2cbMm09mG4Z8v6Vk0YzZ0xZ5DK/4TNXI
CxaIzuvbMYv1X574heh3HHQlSoOI4zRwSKyYutSVLQIYcKnq7kzwy5nypAE48CM2
7De5gajYhTr/hZJ/KacgRT7PylHkrwnz/reeq0augNA7P3mzoe9VaHYb3BYD+wmd
rRLh7AXFkloGSbkzX10t12CdlWyikr2le59LmnnDC13d1lDzy3IIP8vaFcuQMpEq
dGdeMKKFlblHnDp2X0bRdF3T2qZu9Gtq+QpEtzmJwXgsf4xRAgm67KvPzCbqmHTG
3PnyN5+ygjbP9UGUxI3M4pi/lu7Bk75K/Z7rQw5OhxPlMfFtGr+uzkbuzXOLmbNO
v3V2HOi25yQ0k2MdKiRVNu2kjChuV6BnGgecmPZAs4QO251UeBGQ4EeYeyHM6vZK
StRKSFFsC6ozwBIx6GP22axT8z2oRyxD/pN53z0v5u92DYIy8TqTVemd3PakvKxh
T5X18CCSWQaPYgHR4jYvBnV+Dl6e8Jb9eKOejZzeVghs0yVL1tRKZETwS3pYZpWn
upfsM2VYDSna1K5u+Zb9C5BCEQC9GP+szeCQM5vi8LXA113ptqYZaqC1aJVE2TKE
r0Ce8s01bysYb4lvoq+JwYk9VvjNc7kfhl55rVLxRI+VWoi4IbqPbrq4JRokPo4e
vWrUCFKrlKK/TezvUuKGgHCPkqYWcdPpuQvS1lj4KTuVJGxVSUfZaQtrmypac0Ur
xHIWq7pZIjbU3xrCc6O6nLv+/1FYB7mQDO0PKSQoBDfoq8yrr8ZGMO6juJlG/sLB
h4f1b3U8Ordqdxjw6cuSayAxisKCCYtcwcd3VIR47VqHUo4CsZoXRSUBhjjm/pa0
ImdAeT6K+eCTMU6fN/GfSSb90xmekazsR0ortwssjN3M/SSDlIcBPwkx7TBW7VAt
it1QJ25jUfvGn+a9l3JbbvrYGHCXdJL9nL9f2/zY3mWSdkiK+pfMTntNI5Aih48O
d8xxGQjVnEgHlU1ayZZJRk58B9dAdOPtNb79zDOJ/ycRnmsexSmzQhzwztW+RSam
xFAz4HNKSop116DSTWZPshkBs3bRgtzB3OHGlW47eZET2+Woh7PoXSGHv1UkP0wt
QtSAWxFLR/gnEPNXS05Bc8qwLzMTwLe1n79oYuIA7V8oI2uPvb5173YGnphtM7N5
CxB3tWMaeosfOAPhodcm+ceCFnXrsr3t1VaelqjIPUMmwjS5beBABvFw2vDULP0W
l6fxnxkyer5JYpF+RaHYt+doBPkAtbZXTCWRZkNV3sBfOAvekcbvIv6vVDK8TVKv
CXYFh43DC/UIcx7Gewu5vhRDclr2kLVGpLlIP8zs1ARwo0I9ZoYOb1YCh+s3zkAx
feNYp9CY63ts6W0sS+hA+fbBRvjqrckOazl3b86GGVeJ/s56JOOKrfGMwqoIP9db
e/FrcR0F+dg0wOZPJJNyJNDR6phMYfJaojYQeVxsyeoaJdhe+pfarwbqOWhkcah9
lEJzHPkjLyVrnnyzCckw8+erQPTPTulWALoe6uFvO8TDQ3U2v//qJxBZpABrIqSr
i8aUttRApaaU1y+BcBWRHAuj2NjEfkthM5T8/rl5uLdrrr88VdaGLLAJ9Qa3lYkX
Bto/0tfinarW5Yb9aimqIRfb7CGFb49L0XOp8HX27uO5pGtd1aQufYJwx7/4bosY
vPfxIQb1P97GxX1tI7wGrR7AxOdllAxsrW9Oe40125iHHrHbxGAW79G1+l/AnBzQ
9w7ioUnOfVbtrJjxmC0gJ0DHWSqgxDVzCksbS2i9gXtuH8RaH4KO2mDIliA00Myh
pKFhjcsueeMfwJW+Uv4uBE6BCxjAMINEExOPnBRCjfXQhHfT6YkSrfT6ZuX4g6tN
9payhydLGkLVVcGOGGFPBeHUXRQp/E8v0eEMlNMperzJ+e/jV37pYcwd2AfXcjWn
R6ehfHQerDPYMh0RbrWVZs1ujIVN1JumC2dgf41N53+CeWMuDoFcyFAnGPv9dBct
0zCxiZRZoIg75/MfLcNnyeuQhur9bivs1VZETJXKAsPB/H0l26GbDb6ClnbhJaR1
Myo36cy8M0QMyXvhRz4N8/VcR+NhM3HIGSt6a7z38H1cDeACzeaai6GQw+FY9BKE
ysrMnNEGAi9ryvtwLO97MtlwEUB39vt7X97stkx731bUBl9hrmzuNDUMiYJPRArO
fzks9nV0TKeEW1KBsY3VENIBZRw4f2LtXBwZ1ZTBcvkbYgBe01lP3QJ2LOKHUJm2
Xxj7CXyv/TbhGf2+eVyIt8GwNr1SXSsbCmYpgFCcj2qEKioyXLSTCVHjJ68eckK2
3PV1aJkse8fG8kXecorZvaWxGXN2bUSnl/8HB0YCShXTMt0+J6byVn0tD2Q+GLDu
ES1lDN2JPXjV2vFKe71mYOS7s87/pzdu81ooVQkrIPbzcJD+kne8LcE1JGw/qfYC
VsRRm0tAIxZxkKqQvezNpacBEf+rMcQ2XDpNdr23DDTxSWw7shGz8pm52j5iC5vC
sLriW+yGzYbwn3tBM5mndpWUgXG+c9EtQSbqi+0/xPhx1UxFEMNN1ujshJx/tojp
Vh1uUPQ+4kwhcLPDNWgXsQpoW6I2IO+L2tYPHA+ahz/ad7MviEmUn5jBRc0M1rTe
1MRrX6kYRoKYhqns6D3ghjSN+LE77g1tmn2ldkoPL3KKj1AzpfOyfZq10OXX2pZC
I1pFpL4IrW3ZXp3O6I6zfyiVeGTA7VbTAPED8cFzWRHGyt9ngmJkRYs3F+7qytmV
OCkK/LMNeXRZ7gfBquM7nrIZ2EtNCxYMAYyn/v/SEk7g7jBwmBwJwrq0MneS4LOb
EkwiPRqvA1Qi1pgzRuTXUu+c/8JJeHuwckXmX7Jw4YovRC1GaIWdJZtzb2o4wwgY
yl/9djTB+jJmefWNFl2ijJUfYOCGwwXdGO7IWe1/dCiX3VfXAnL043n6q/+Pwj38
PmQ0EQNcZjkTRiQdFPJ82ZjmLDH+xfj7grJGnMFSnal9IKuNxgDC3mBUL/OL6krB
x8NxlBO4ZpDwsQGlG8egXPJZZHoXsNRGmfsHL4uRuInGWP8Ez3Jzko8CdDGK+akF
h9fOlqwSfbVFSIDcYwjoKamVO2igNSGZ/OyywqH2l/07kgT9+iMsprrg7dsifEBk
e7et11zPeX5eLPYE5SSU+pYOWfaiqVUDIsmD4cDe/w8Ib9yTO6bwGM0uKVzCFH5y
ual9Bn5kkDTmFfTFxCEXm5xDOaGdSoP8iC65VkFObni1KhRORCwV47rqqC338Uvy
yHvBn4Ls+ED53A9kQj9Hne15P0kkdilMINz9tIP1EEV6hplY4yKbGi8at/uGwrjF
Bl5TMwjf9Kb+UqgNBboYq/p5XN1J6DiBVvrYPyoI8ejqX3v+v8hMlWPZ0lLBsZ1m
LiDOZd+c50CircyEtH9O1LHpDJDcXsVIxTryPxh5nUbFbmP20l7KLDwZ0DvHL+t1
T/nmWlfs2MKh2HZ8MrCtPl+mC6lyL6DBEcxqF/WJDfPu/DZT00bU01xyIpyaHCrT
JvjGyomn24qmJnPqpLn0yvIyBoAjlS9BOWUCQgVPrGm0396BR0so2xvb4qWP5a55
bctFXn6nznVvcQrdkFT/HIZqzd4TENLsy9Ilb1mfTIQGfSXo2v/5xWNdeSIkjrXJ
N4V+WzKJ0xkzllT3CI3c/0APAGOUe8SPBWiFEo6iy6a+ZRzdGE7cR6V/pLFHU0sC
iIugeDNc0PQ2lOZoWG4Qr2dcDQA+uymyRRUWX3Q39oe1yFX+GUwZsS3+EiXqePfH
VLhaYrHNIvQb1jOJNo1EeKg6RHGt1mRuUQrZT7Mno4i39BpIhUDyek9oWQt6b8Jd
0GrrEYd3lYTDYqcBMFLrQbg6ARKeTEqHMBS2sLy4c+ElrK5M8qM70gv2y/w5pE8/
vQDCqyYG2/G1lUs8UiD4oW8aLXwj9rBZ96SF0/G05QRlDEaEpW9+TsCY0Y1f5tu9
/cTpGhkzGABuIWxLeGUhhn8tw9eBuXQ/rpTF6CGxargnAiTXr+vakry6k11gGKn3
nlcq7r32dYrvBm312HYONf22zxq/b3gFPZpxS5albgVW6/963gNs4sBsKmJRkMIF
G17Z1oqc821HTCwfkuKnGAKib0cOZv8vFsnAHWkmrgv32qvFdLUggVH+mALZ6HnA
JSeB29CEc9m3vNNbJJqtgiQADMYj1QkPUQnEXwEniCBhek5fucfJoHGrNKnUq7q/
e33KLhU+/HO/LmUZLNQb1n2RCBAX7U6hgjXB4T9PnP52Xbj5xuhk9nF6kX8Oe6PR
JW+quGEhu+Nsz1SXuJxTlnBFtg5tkzujUrl5UmWivup9ff/8or/f185IFnr+V6YD
9TmGqEB8Pd23lqu592yjE0EYDGijsQDjBbp2lbGcEKSy1oCXz4R92qF8nxFMFr0c
W4zmNZjMJC2BRX87VfGbVG8LiZ0NwB18HtQIhpmojg+hQVAf9Tn7bE5UB111cKSD
7ws2eI9VjrVuN1UFmqUffAM7I7YbtPsgkE47DwBTV+Li5rdQfE2UPpsSL3Cg16Dx
aGlFWjvEWt4m2JqK3xnA2htj9znbCk2bvpbJvv1n0P18quav74E4bJHs8eLXEKEl
E2/Q/Q5AnZlWLMxzJFRBnIioPjJf1zpiivPBxQWfSls+PtfCmZ5oQ6soQwGKFNbP
ScGmCQw5y2u2Y37CbVwcl2xRJs892xOkDv1iF6817pvrBOiJKREpRBP4Vfu0yU7r
hi+idwfdSi1O7EtngJlsvgrdtDBGsWATWzB+TaeOnmxx50k5O3wlGpljOwYsYE3o
eiCII3NwIqdREFVJff7iBztYpltnEXumnCrWdiIOYQeO39eHuftom4+yYpqy7Mwa
c4Xge0/rejTRw19HkHZH2/Oyn3zuzV1Qiv8aEF7dHHQTZLv+7ERq3pXWPw8KUtXP
Hxg9t3PL6J3cBJ8oLgODzJVM9mHOt6dqwH+3ZT8rcn1SkPVDxeblG7Z0+Ad5zgd2
V86cr0EgeM034My6TNzlBnuodNtjLuqTiUFBWzhZb4P08qgGFynAqYGrqEQSL5il
M4TMOdUjYJYTyjeEKFGkRyNXY3OmycHlK3hnTbs6ZOZjMqKHE6FDtPPq5mwh6bh9
npS2HuRUUgm19qdWAIL9ogPV3iKi/JX8u6c4wGxb7/p8eYyf1lxESd7VoKhTaikK
WislilHOqGlkhp2BMYXD7/WO85ZG+ujp4D4qJNPoOsab7fA5uK1sdu+yX+c0ALd9
wtmQgXYeS1obW600fY/wK6epdAFYjJW0jiwREchV3k5Uaz42QnZ5X++1nt51XUrq
LgDyPYDsvzPh+fnDnzfZ7VjOwMgVRsmR0Uo30hxeLAhCixchXQ/FNbzkQI/fVCZu
1bQJ8qVzQGBrgp4BT6cxFpOw8Ptrc57yJ3eenKrfgPcWunnXqH9JGmomJgRdyj3A
V6485HX5I1T9Fb6F8dH+TDS0MnfgHPhSXu6Ou3C+cEm3x0ODUvmmOtCh73AtkJrP
qm61F2VPu3lIJL1eiQ5Jpax+nVwiogZhqTJEcZ5E+AM9XZpHXwTu94xcqSX4BCmR
ETXgI6u43mloW0XZlwSBrAY29a4sesE/tAFjkFrw0sGbGoiWRcfruAOAKspSAEow
y9/+V8IFnSyj3WMWrXLb9TtL5o1xyPArl95i9e6eVziNrDK7eok7XOlZhZAI0Frx
YBYFpnRBmTKpr+MzLbNrvV/PsN+a6/pQJ7awFELrRR2iGLaZ0b7R1Kl0J/84Iyd3
CqArTxyCa2WPjhErsoy1QLJoDXiYqAMvqOGU1R0Nx3buZMh37I8z862DLMs0sWPO
oXMzr+POVw/huD9o38crRbuWhlGb73+uIAiRLyAhMz4f3KsZ888DQ7ENtdb9yNmk
z8q4S52wN9bhfkkgIksV9gQ2AbmbBR9aVCOc7sZRYAoD7qP3KiF+hbtg81dgY6G+
G0rBuwavIMU/mSzHIHLDazCm/xaWeEEHVl0sJLLWBbf5PPR00HdLDtrSBf2clpyf
+G9S4s4MSxMpphvKFmq4NERcy3NRI8y++DLSwVk9TyXqj4wtIp1BfTzCIAnhLTh0
4VmVI4l288jrXfAvqFVbZvkwE+ex+t1dR2L/cudYHXvyoQ8a0LksTKN+HzIPpuIG
NDyBVbJte2HKZhnaAK/7V3y32gjqb95Qu1mNX2Gy5oTzjyCz2k+BHqWDID4G01b1
1DQ3xIS5fXTt7oMrkM10tRTnk3/Fho+Y7p4WlwXebhhbQ+c9RG6Lo/XorZ3UBnRd
EuuuTQbCsrwXFh5j6uSF8LWVxm7wmSFJce7xQeSCzrUliYWWGahj5t7FFqHpYCaZ
GrfaHLcb6Plk3JVPanFAx11Qio7jfeIgPjwvRp5p1vXy6F+phoTM/gxA9fGN7WOe
SgHNIJtICkoF88ZDPPhMRUScMbokqdGbBqwK8GOuqQA4TfbyoJZ/rU0ovQY9YOzZ
xgZ4bD3PM0yv8njT9/h7HfdBjh7VMtSIS1O3ipgHZmNM5b5bBeFSO/T+4hUjhPfL
YqX4uigeXGrEhb4aYdsdOKfOo3LDapscKsGmsvSWDywpZkMvxXDKMHmb8Xf2N+iA
+WYrPXKX2VpVABdwEJCy1UrY6lCUfUuef8k2Cv5zgFOuFHZmg9hg3aOmrDVKrEuJ
0jmB5mWBJnLSE3pKlXt5dtjNKCfzSYDKTsv3GwWSkBsD1oFXArXdpb7qAGvFhId9
55ZLO3Yt9D7zORDWcpWbwaTHF1jpQcGTe6fT8iQuvf4Phpde1GOFnCVNxrryHogj
YGL+2k5lt22aHmMpGxfGSsdbHXtE3w3ypsjHvJiRB64j1zaH7+eQbXu62flQsbH8
UfmlKYZeREeN0AohUC5bOi0LGFHbpl2e+8xFomcF5xEoVg4Bk78zGqC3YEAHJQNd
fxtMaHExHAIuygQBHP79D6qkm7XM5kxid4bzTuDa8iu49yF6qU34iBx6EQpBhZhY
loe2/AUumFSRirv68m3pw3/80RbfNfXDVvaLrWKd15xm5XvFEWVExV8PWSByf98q
PwXVyLFLNF8qQqeF3M8GRpWW70YTIhGZVmjgo832/Oq3HcnCrS0Ee9BGIVqdld0M
X4lAsuE7QiuwJQqZ/TCkRLTUpZ+skSb3oyCH5poZzZAHsjUCphbQ2vprp98OxrA8
1Yyh5HIdn+TBJeeP7BQLufWbIEXKpj6xdYyqiu1s2gvSvUvGSv/bVxmo2PEuNN+u
bMsS24UEaNeGuhLI5YHnccLR++JsJzVylLPPl5htEf1kqfdZ1dxXxwnZdziKveNz
aL34ptyli1QAdS9IFm+5O1Zd+X6L4bY16jThA+pqVxj07HR69C3ES4flKpSYD/kE
jvjXA4uNuYXMJhKM0cSI/TuKIt87nu5tces0Y0G5RaC/VWfQJ06scc/LJ8dwtv/C
BEt2PPkqIMyGDRlannVGXrjp2sjvEgCUjBNzcP5bAhnWEqhBFLewxHezV2S5utN6
GYsPsl9ztt6sRszl77Uej4o//xfHp+kz//2XLFOfDrO1+JJl0WzFUZxvjcXkqfhJ
6tdoE43X+yqV0IMGo3z5bL8uzTumZQQguHjLdJ2hgLT3XKY3d1oGJhzlh+yElOtg
16083pYTIJR0JViHC+KUNmGGu64A9cAkpCNpftg6ee01C5K6B2spCo3va263Nra0
xZyHO9NvhRfYGewRVKHYkf1F6KnmYZJt2fN61/Vf90HEgwtf+pe0jFCC3r/n77jC
+afycowXogi/MhdToxYAMCsQwU/MhCAlgmX3mKtoYc1Gz46X9FpJ8/BFZoZX6jGP
JP060F4mJPrrZ9q9c8rO64zbkHx+p3el33j7vMvakYEPdhdLJAfqD4RgY8jn2ui/
E6hT9Ch+8ExWHU8Fgeh3kYwbXfeLGcrjhYEjvPvdhKCveF/JvV62O3xA/gEX1fo2
CRF4WghHpZJXrieE1aT5ORbpvLJ9f73YZN+8lNCurSLxcPoSgOvb4BTVJbYNYCig
HuwL+EqaKPFbEYNyZddgqqcCZTPl7C1EjLPc5G6HyE8x3epyEbETSCqb9VZMFKfk
AbDmytJG2Y/qBgfHhC53CDwv4M+t93kYqyN3XmIs8pMi/nxsmq1KLaNh96CF738j
gc5LCzq0uPLnN9tjNQwg8Hr+72z8Aikp6Z5+DVa9swwy7/eF+db+dNw1TKOPaLpS
6M8jWjb+Ah4Zrl4dnzN2WT+GYFoZYdFQR2bUaKBZUMoumvsX9oRPmxAxcOmuzrna
2nS/A8SAp4sQLbDALn07h2F9knzD3MmqunjW9lUU6QCbrZWDTJgtcDy/C9Q9BMQn
ADvYzVH7/KpUfmhTyTCWJ8u83xNCWMiNyH3kt5sN4uFIxXAX6n3Xv7IO/G4QjNte
syPNXzOzDAnen6pBvMxbfZe6VK1lj3H+dVjUX4HVjLuHbkT2C9v0lZx7h1etlUfN
NNeZTDeMaRGhD860gQ1mR6DPjSG76wMCGW6HergjwmULyKMOssOom0Z+wEbb0tVs
msI0mw/ze2AD7E6tbtLpMs8/6ohuBk/eFjoN6DLj3ZPk0UA1cMYV7JDhbVbnaycm
RbZ7pmaAVEcOFA0jOMAXMwg2mEwdUb2It2cMGGDV2J6rgmSj9O5s44kwisii/+GZ
oEKMlYU3zW+1/38iDYJxd9xfisJr8H3PxWVQjbV5dAwwPCIFdzcrgCcjh4DpE9a0
acW/+y6bpD9GtJ9n/CDhdGcRNc8MTb69rg/QbL9A2Yz3cEWygTVLgaxTHS5w97R+
RPI6kBVFsBvixOYaQELxGVVMZZuemIffsf/zH941lDQBRQXPbakyAQJJqIi4cJSv
PmKUp+jUfGD3/xzVxMxqQIHN4BCaA8pASeWRcmAPb8j29ONEG0Z9CIsaVJyz03D3
OX1bNtWcF0W0jTpneoTugTz7/112w5f8BWT31Tc38O3KdqosbFgJMnSdpaiLjbLP
kidrdg5oK2wtOt7iH7mNySI8lhI8cQ23qwkiArp/LjopkU61k1tcYgQSfMIcfa7Z
5uiwlfNaO8KzP7V5FsIfhbpRmX7Xzy4p06bhq/VqPrX8C6sbKqefIyo7hgC075sX
Q7AC+CH56ODCjVIilYN8COnOUoltZ1NZE/UCy8s92XB24s+IVmp2BFvimDx2s6vt
0xipZzw4VLfxhfSGGiOw2tZic8CD8u6K7AtOAwDQSG5rV5bc7G3fzKuc8EO8hLr3
HAEejy9kZN8X8hJd1+MADnug33ijCyMDBGh2JmxO/uLROqeT9TkWVdO0KGS7v1yN
PIY4qQlE4EfFMKwzAvNWKu/DkabScPo+Qazk6gfkv/fG2nGTVTjtjublUZmu1kkF
8UAsdvSFswexlgJaakR7o50l3S2NhBufUcrhL6Ox4+1n4gFGuXiVdg1ObcNb7tB0
7XI0lQrOZy7D+mU3iitPUU9+6Ye6FQ3p9Sb39I3M0PDwzUGxh7LPuM2BS3PCNdnD
DHSnkO5tBwi5ThrZFdcBBOG5M59kwTt1wQssaSmJhK27dFulQP9N/pgi2LyjygJ0
+YfmsZctb7c7AOTnD8ZPZjb3q0ba0dTjXHoLfJakZ4pvE7aah+PqIE3iwznL3oyb
Uggt51pOS+5jUtVqKx1shM2HWaQZzrsWtQJCR93umw2mSbvZFfSlwzhFlmqc7GBV
kXE1kfS4k7BxrrRzveY1U9EaijUNcr7QeSbwquPtjKmW/XBJrb9XyJQP4tr24V5P
fQD4j1r9vsKU5kUqhTu0eaMoudeHaLKbf79K/xV/45bWP4xmaMKWTEFz16Q1rox5
ptn08J0HBABHeYrDzR46mQp/S/6o6GQAF6HJF4MXK9vZxo6LsofBMsTLZO8Rd+BI
NawVzyiutsmv5fOP6AwtKGjNr3cZAjF5kMdX5Wrz1bSjs9adTpwf8J6f2flQ3KsF
QF/bocrV5lZDEBnwb4RAic0bJWCTpuP1EhNrFenzUDlxX9u8DlMZ1tjMTi4bsh/j
W9YqMB8qkZpn1P5m2+XsWJAxQvBXz4WFhY3oSjbbt3J5JUuNdZpD6VZ5PTuGHbfX
Mf2FzmXQBF8LOZmHaugUZAxqYa8goBv5fQRt0kn066Q1gwWh9i4RhtYdJMlS9YiA
WUChuOW07VcPEHp72UNyNKIsh47MHmR3kP0NnIL8MCn8MhiIbJCJ44bsCoivTmwz
J/RXf1Nh5rqL9OVTfATa9mr1rGLPhqvW1ZtLIUBFuvxCsnG9AOQztz+bSJCBExcZ
JKqe4L7RZY2zZ1hQXoArx7uVwxQIFLhY53kT9UEuoTlgVYgHUbY6Vn9/0fVqUdMM
uI5gSG6M7RaTYzv/MMw6AkJOnx4a2lIYKQxsIsGkV0QUqe4yFqZM4+2sSbNFqSVP
Vmu0mnAZcks4LjjafQulIb6J6gdLv8EBTo4rafEnJ8iMjksXCTwBgKbh42uwDCyb
a8lwdDtMLkJ+7ucU2ghM/EZiw97L8APH6dPzuCqw6/wNsUYZ6o6cDdKMuKDSwm6C
fP2hoQV7D7FnIjZZeUCD4gGL5c4kC8FYI0RV6+fijfW728WaNSBAdhIH8dW5mU2l
3CqFTnX4Gpj27979x8EuXtv0TZbWcTBMHo/+9FIDKfKtSXySBA01V90CwmRsMM0F
U5u9kgs1G1B936W4S5YDSSrZd2giOCBS/BBd9X7Jo2qcsWCaVl6TXo5rCrXAAeAs
2MgMb8ARWrw5SBzRSk3VN+DlXslsauvQ0jiIT3sJCOLgD0qdIqO0dBqf+z3fREfL
ShZ5x5r50V7MvXemZgxgC8HK9WRaUmA9gmT/2E+QNwuMM27k7B4DwzdrY55SBgpP
X669aqeJ/t75oOuadKVTDcNq6Rr6daoaWjB8zr+qszkeJJhVibPUvbKMwUjcGZa0
ZkUfSnlLYwUek3UTaFfQM6pQCyVHuBd/slAlYRfLX0MOsifRSWa0dZdOf3geqWzc
Z7zDbSy+ABs27eB7D+GJJ3NiAw7uYOgY/6K53wMxvDOjLmIK4vR8vEDlsKS6vNRH
POWsnlWt7E6+frbIXPsDulkZRCbSamc4TeFesmqt0CfdO074FGkBEZTjZHRRm7hU
gFgLZSDK2UJ2EJxFtJ67UNIKmqlbXXXjj4GW9VkIrWaMtJSiNdLSNKa+755vH8gb
GCE+a5zetHjNxLFmIVcLj4toIiDeOnsm/MMX+uJ3aY+xVoVHvMqiOSxTmezGqY10
/08FX9DxbxHmFCDUzJapW+X2tZtHVp4JjW5k79muA3Mm5q9HHfbAkLa8JV1YPHWf
xlHt18gImLaDPjXOmIn6yR15ZH2wWrCKjkht4UAvIOiWEc5eR01xNbt+LLGKMCdG
rszWqhTFvXYD2TgIX1p1/iyFqRVSkoAKe40x2i55/IxvPveAn4tcBdgz7XS/Qg/c
j9JRiFt2NdbtjyojwgC0W3BETJBUCPE2iTC6mX7yS6r5NhYJtSWu0mQxeUHbMLrM
tcMzqybRqTh3fPD0WxXGp75eleoKYWIrNJM88t8PF69aSKiyEf8hb0xiNT+i4rz0
IQ7ScKf9bYEvuv14TE4fyJIos5hgckeOhsnAwEmBnDWJV1fL/oHxPFFsLch925pK
IJL1s9C7AjNJJ18Cd0UCqe2npCuNXqq9Fzl7UieOta6yzWXf/W88lDwIHKuk90MJ
Oz9YMmpuaInkbgfFAH7QXP9QFzcb4kIw8Q5hhCxRzFBiEPSfP7QUkpcrMKVV+gZv
aAZwtXxkQY5eQfIjCNTMivfA05GmtQnBZZk9R09xIW/KocPrd/EBKKVvb1YYttla
5HoPxVFX5A40oNh1dpJps0Ky4x8rUs7Fii+F8O0RAVaVAjNExSp+iIFsqiZ9Stc0
+cfdSK16EPRNrDeb310ak8qdHcs55eYGKoNFzyPXA4320s2Dl7q1DgLgUxS2u0Tt
KewGDsaO3nqK7hyKGnCWHiDgas67doxMv7esnT6gsTaPLsGDSAPAUZVqW56Ddlt6
WhNgqhRAlIsqQhztZICJBtBUgb2lyfnTbL87e1M3NC/1yaKCIuTeXhR+4yOgNJcf
xOckZIUqWvWnfxRzR4JjR4vkjEoRZ9nPwRgQDA+yrpkLl67aRWMY7ZiK/QEzDPE0
1Dvjn/ack4iquoWMNyljdwd06WVRF4+gTGOmB4lIOhD9ICgojNYikB4CZ3dvIXpb
G4JTC0+UzNqXF8WRNEFPR2iwopBg6pBe4Weh7MOf/SJBy4consitevpiKRZzpgFi
T60ApWolDgSDIz74fMA9Fzv4bw6TtUPDtaC2hkg0Q7nMcg0jRXk8uigE8CoUmKmV
o9f0fLvHd+AF4oBqjBWI6Ldh7OEdnBH4b/0q7k1p1vq/WNsUtpGr0661uofvyAWV
KnevAXD1ASWa9U0R+BLSrwwBNBmgkJcMFllOKPCFxEvvZLlLY3D45x47CGXCMFF3
ssxYk6g4mTwS3ygrYzYzqzpJ30Xg+Pmn2OfKPc+3dVGRS98fBSYw82um1YZTS8UF
dI0sxra3rK5RblethBTljgSX2W5q/K3bA7Ho18BgXYmcfqCcbxX+Z+dKNzURO8YT
otT4YHth4682S0HRIexdR8n+0h8KUT6RBVQa/FsMT4Z2IxPacHZTeWWF5uX3DnK8
1BfUxLz00KRpxKzJejzts6P+UmTJaK0IlIr5J7FOVu4zFuI5mrD8JKNAvhT4J7Qa
rftX+7qq23as4xAls7Ohcq2ZUPwGr8tmoAXg4q4DC4F/Ke7BJDZ43vvkW99fkslB
PDEQkphc1HYK71pfD5XZopGq+kROc6Tf8k4xy4Wj8QPxPrT7uuYCrHptqPbT9Hsg
gQij8cf3lPasjOoTjTzbh0LEgrNX0JCtpEIyaZWDDglCxyUWIgXUYZ9cReMtbfd4
33/rjnSPoWjPUiKuM5kOrrP556zRiyq4QcclKhuPLGyFeJwcZnnJjk3DDDnk3wfz
LcDDPCO7tMee0hx/y6C2t8/Nte7Ut9JToI9bbv8T+QIHoW9aCGt/LCL/Yh3QXEIJ
BtIPQWLHU4EoAlMhXwsaZOoHfRsx3Z++lFqnbCYegf9eGzWXjgqpxUjhmb8gcmMD
KdqKl52UipYMpHVfDIu2TUJ5klM3nnUwzSFg0RX4Yc8z2/hs61A1Lx2XKNOty4NZ
CG9fl2nAIzaQARFS6lsJ/Y4nDUuIjO7LHF+RADqM0RhVjh3LXWTCFsqH7RL5MAOC
uB/pTWtNiUWEXCBDaat/bt2XESI+Xu3tqRGLEYTTIPG5KZ9NQFCW+FjajXkuFXmw
ihbC13Fi5RWAk+7Himbqf6wcMsiPx2YTDCu98c/0gviDKU1HyAay++TaPWULugIC
ZRqANBqc8du9bGsVYF7xdktGhkdk1WHV8uukFvgaBO2tYaVEu+G4FaH7ml0kVHDy
6bxq7hWt25TvrzEtgrwq0v4nrUi0QMadZ7fVt/JmudFjuHg5c5fs61rfKgRd57cJ
o0t5BZ4xIAd6CgQvTZypL0WDaBlgGJL3wjreBRGyBxZvEkkTgjxBb4iF+cNBSZq9
umj5dm2n1zzwMGqriwCOnV9yoPHfQcCqHUF26J66SF7EZaaO2GMAozivlQi4JTpF
XXz5XorFtjGm3a4PXtb5JCL49CfM2biwgE4Lr+FIjcow/hYHr3dFmLrM4B86TySh
QLVOgWVpBiMSNmi1YUX6Zylns4Ne+glZdR2MRvcsRnNAJSA69hHmJMVOtj/sH/jh
fKWYDUOlHmyjWZ5fmUix3Q2iU1sXCdwEBbbfpzZ6rodSABTgUHP7YQmp356kT6oJ
pw6bvs3KWhAqU8wK1PH9szlScQih60jNKqrRxvuN5bQwU8Imrqf45kT2kivbOfdl
03hP5rAnXxt2nopr6+uIk+ZPgTJoORlQo7AXYts9NbRiVfabzh5dYk1ZPJqNOR29
e1YDnh4ekaPzfgYjRB2J33dDme88CGGluczlwsqd+88BUqA+SYLc0t2XuQGoPiYP
gt3+dIgsCLWQLrG0k3BuaHSyVzuIuL6JpflUYR9ZAvFPus7f4lAv1n7f0+OoUOy5
Jm5s9/hbalARRimCwlmEElvF/vhcdo7VlsGJyXrpFZAn9ERqYpfWehxrqThOhKvM
/i4Ev++DBUNaBUcDZRBdXeyaHi8SGFuBKl0srCp84xqljiCQN+OitWagB12EZ24x
DbY6hkEWIpqo2afGq09qpDWeXWa164goWHcgDHtUyTgJ83g/8tCDYzMY6YTCipEq
bXjpZXWoeKdLjrRYlLFJzq3QK/V3BQyPBBo21Tejnrzk0m5ZWtPn5YbCNaZfWopn
MCblPPX3Re9QHnOHeKhnhLX6ydWCGOV4gb5XHcG5a7zNsZG0lkeT8MDzELgbmGet
phs2lZMiQGhjE4Si+4P/h7D+WSt1AulzOpbhUS5mU8vG58+mZeAKyyMDgqM6dMw1
eqTaAiniUywvgCqOaaQORGWjbZvz4BZuoWGggYdt7oHHFIcL19Zho15HqQhxPQ9c
Y+TGJGqgwe0i7S3Fl0IYUHfEvRIxArM+2sPSUriyBq7FWHf9o+zl5isQEord35wC
K4Ky1WlGLc8WKe5b+LLU6+nQhCLzjhmJfnqgROdGaYPSPvx3/p0jL9Zd+2RdpEKT
RxNEySheLieWo3WASM19xAGCjZ6j2vSvt3myCzxuwdqCDrZkvbXkoYXEvhOynJp/
3UF/hhd8TsOt+OXOtn1WSszFeGXWLsVnsxLZk0gRkcR91qbbUdTDOMk8cMZWn56q
s+opKUV11SZYS52bsMiHNlo+Vbohvb6/c+VmdVqvTaHx/tO3p1Nd8yhYANSrLuMF
hjA9eWdO5HHYzc2kA0b7zA8ZtHVcduA6wMYi2NenZcRNDprv1ZRAn6iWEiLtdVIy
magdU0z0CMdLXltJvOYCLzaz02rJGHIjMoZcemEnOasE8Qb3lgkw6ksVzOvjNT06
wn3Hj1Iz3b3T5Sd2wa1nEpXHaed1jh/MZevmC1mbAm22xy/9iJtUg1bBupnVbVJX
IkmA0AqVbQIbB7fbtiTFLDNc9WL6lbUTPkJGbwV18RcN8MWR4NsnxYW9oHEqD+D7
ZhCoeoLvYenW4oVmOajx9wwpafVZ0W4+q8iNgYHALZkzkCedR96ylradOJZwdDI8
xx3uoEFZeKonR8cUNRM5PH/ETbG6jHdp6WVgKScCIBS72Xi9aNVuib4y4Mmz4zTO
/cczQMvquW1fBIrmg0EYFiFPPNgQLkoaHkjvsdkvjtFa4o/IuAnHdEqPQYcQ+3Kr
NACdX2h2KCfThGSQZiN/SBp2QyHQOVa365d1tf5abWTvHWSG3v85hqKTMF+pumHX
wUyiHwK1/IPTS8pbhKp/xa14918/oX65EyqQJgUAH/V1xyQUrqa2YlCYLRSfTC6k
lAgw6iY7LHstvssWplrvnZGgVy/rM5YAQ1nkfAceBXqyL0WwgboY3+y545FP4peA
FiHvLORNcgYHLLgpxYyyTPRoo1f5PRFE1tChK87rqMa5AmVLX2fMQdtRQEbErGEX
d1qph0kkeWTWIASi0UZPPpRH+tVT5L9fcVk9pkt0Laj1hWrUmHiUGOrTlEZFtLH7
d3JY7qrCzumyEdzypWO9RkFeDDfAt39uVbmFSO234M52ZbWIDt/CD6Wm5hbMurdy
izSFOO7rsqCItKyw/tfhVfzaeHe7E+Qn3QhlkBKNbWv+rcgAGemgQgbIq1TH7fop
wZvhEYFwObGdtyMCU/0zi6HUxz0E0BKsUnzrZuf/T38RyAYOeg+hLLrTTAOhJ4AX
5maXnsxcpiWAXs/zWKpso/GctjUzDcC9mr8JHaFnMSrCNvuns3hWHNPzKPqonwjU
P1exZ1admMtq1MVs1BuCD6K6Bsg5asCiyNFHr5ndpg3my01lWEiZbidSgEekO8BZ
Ztm7OSLSDnHmFJY1Lrk4RD/Hj+fRaNtymzbulb5bNnvGa6BQkbVsdnH+txfkHbxY
vkhJCHmh50ruY92c72QecD2DstE+A3wHacSA8sddnIi39ZXMxnqiVFS6c7UjvOF4
VhwwSX9zNOZIbjHRao8FSbXztQts1kpB3e5UIKF+pLv8RDP6tnz0YNoB9gohl7Z7
MYSmgPWL6YhYuZTSsO6S31bACN48Wp3yuFQO16mGYAquhNRba6LvRDmtKNPVHpwp
3RIq8nVT4sF+fTt8VhLuIJ1HRxAYvpC1QDAx5sujSoQSPJ611JfaKj/E+bk/LTQK
+QB2ba7iIp83AJrJXmvDOpwYisVRv40VjZ8EhgnnzLOAMOsuoha9XIN/8XWZGRIx
G5zMlgSnKNu7a13cpWY9Sl5j6EHpW9Fsrf9AQQmaoyxetWgPNTgJuLAM4Zh/flRa
Y7Qoh9z6kQ3MxoYQkCg6oRXgMVJhw0NTP5bOzUI4dPTVYwyaT2AXx3smZ/LEoCA8
6w20ylnMsR/XQyEVBs944PaKe8LklOrlZGE/bcYz+CDahh9Br65uo42RFqx7ZFzS
OTqodTddItuUgf6wwUQ53qBMpqcvxVcULXvyr03hrY24YHmfIQLiUmaPMF4Rdtiw
4UbRcnUqfnRtV5OETXyOV1r1W6nP/5eXEyhD/4OKaYSVG8YBRFmwK5x1ntRUMrS8
1tlXRSRj8OSIzuFNTImaErKC+cZxGffnXCQuxX9U3ul1D0ycCnuu5NN0OcvJHX1u
TH/ZebV0rO5jMRAgPeGmtnXXd8+CNUdDJdqKULetkhkMr8UGZzecoAHw4eTE1Dso
vgSd5FdZpmFmzGsfBwLhcKuR27HuK/oMhTCpwqf+8E1znVwIY6ENp5LRBcc7JqX5
pu3qIjg4h8AR6ukpeiVml8lWprKGSb4yfmSY+ZwOenGHHRIsC+whSB/KezBWMP+b
6OZaVLfd6siGCT8wisqlABrzUOeceGcr5LzQxssIp7tu/pULTlpWP41QIIkMhenm
7HHPuJIgRECXjAUxbTyxwKt5TSXhHMIgFe9IW+LWwgf5IkaLNpehcGCP2JlaaMDI
SaoXltlL04j64dqTbNx/np4RPO6l1M48yw+JJS+ouGbdcOAhlSpnAJGpuRHx1nXT
X88LDBDFW2SXd2CsgJ/TPCMrKleCSa5qksuExywbU1HVLTd7cI+kZzX0JKd/v6ly
ZSoygxArs5UoxomYj7pn7tbxIBRjW8j/G71A8HAfchr+dPo3oh089D9NM+ZsG1rX
FLzbHpYpNhJAkGQ99IKY7TddYpCzNKGe8AoisFwL3ornH6CR99TSM4DYUe8cvs4J
iNCXDBIlMkUBuSD1vL6jrYzDFJ/FUX5hIxgnGxDqmq8AOmsW9fSQIVAleCcxxn6w
7OcDatt2EtduMw2Bdz+YkuNeyVCEDy+isBcQz4RC0KXohLXsATt4266M8dxnHNnp
6aUHxO0MF1jV9kHfCa8eg5AhiD+nBGKONpgaS+28lltS7sxr/gYOl2ztOW5vHRFF
BfwLQhGoIUUCE8zVCz9NE8ALotvJtAt8v0wgvHiLKcFOizddxQ/M37RJnxPWZpkv
/wpvjsf8OikqBCyDrYuqRMIIvgvcv9kOYyni9r08JdGs1PGAX7ZMkzUCKuMSqRjm
WOjAo2WpxmrAynkz61RSKJ35fEiE5C9fhGUHRC/eXxZCBtpJjiMISaMV9CvGysOc
7vHpx4d6a9F+E+rHApmvaqMHHwU6vXZARlxzW4Bc3hOirm2OWrhqn88OKVDUW4j2
4SApVqOCM0oKI5Pr12OJbrUqGw7ifquRiwuSqc31xFT5pKiz/BxFPiG81yk/kn0i
s3HgLjEhQHEBF2kJHaxEA32n7BiT9ZM4fjh3kYKmqwHwCoRpQ2XcIqhGTgfiod7Q
QJID5FSaVhzaCyDbbAdXzPJxHu0rtozBJwaDeqvYC2Qoy11AJBr1VWMG+C2ITfJt
5ZBRjxNzx7nxXMi1NbMIWZMZoKhBec6BIBQ5OTe9tfH/lnoMAw6ZkDOOJZU33Aue
KQcuyoHLixIQiioUT2kKT17+LvDMKTTF3IrBXdJEZxUABFGkT8jGLn/QkX7LdKow
7CEALIxD6xg9PBMcPUQ4XxrEYCbEIHvQMTjQ1ifV3JVc7xph2WsDtCbZTLdsbzXE
na8y1YHKZDDdRPq4wE9ixVSTNcGDXUV4pVNimAlwa1Omh/iTcK9m1IkCLsP+fGVA
OWY8nHnrx7tUAJD5w1Bj8/zFHGBnwcxk+a4bUTm74w4iuYl9ZktTLdFJepxUDeq2
jJr9rw5sOJ3MJG+eRwjODAYvLSLDesu/U0jeI7bwApFzS2jKZehTDtDSGXWhehNQ
HV0mAmPzq9V8KPGoSaeIRubdI3H3vtemlT4UW3Buc43H9PelUvk4UM+W4WBtzQWU
TzZosxfqfbbnvzLA++vdeO86rZZ3GQWMhrnoU4STfrgDpAHUNMqOwAT3OhjymAV8
YuLeXOn/irSnCfRl2E8xkEwY6bgGdxfTbUCPaKAwbjZ7+bMXVlOzAvD2F7SrE6/f
SIfEyrGKQ/tEHHaG354xAucIC0CE+DBQhr/VOJ5QO/fhcbpFEtLKY6sGfunoW74U
NkBh+IBxpgpUy/wa8cvYgKl4kTkICL/9Vhll639LtSta66RDNq4CjrzY304JUcAz
GaRsNpiy7V8gD/Dz2iwmM9bSUQamBGuukvNFGRFDRBkOPmBt8VIMvtl5m1j7vk/r
mGRpj7ZbLlOIojTRL56rY8PD0xpAsGk2PCKwqHvR+mcxaWyyJM2AvxoHUuK8pmEl
bM6W41StwnqjnSsayjURYG7xttpv+K8bLLhmZFW2j8caZDDExXRe3Wbec3CzKAkr
Emh+UasBhFGEKWclxxi7YMs64uj+e4lhDmy7C123QKGMPMQyWTSxq27gm2YaPaEM
VaKWG3LE29YAhTmomLgjJ7HQjlYzdCrQH8FSYbOR25WDjXpNJgrrmnGfpKOPVew9
MzFzEMEgIC3jNhAe0OR2MLSaAlKtuVHzdqmaEe/aboVQFN7dKbld0XdtgnLH8Z5P
XEnwGZxCrRKppi2lK6z6DsxpKMspyBCZNCPbdK0+1XjiawRSIqeZQ3btwPpOYEhi
lI2FwrnjyTFct3udY+bI2KO+fGBJF2Z9kTn2DOFi375TLWdxPl5SYtpmX8hFcjx7
L6OK0iHO7RsWUJWSLCByq0NWUsQ8DG+svewgfXcAjYQ27rOOK/5WcrJ31v/90R7I
1kapvEEOQOeIVXHOkVLQv0Lo+NrM0BT2cIbh48UbymyEQYNI2bIvjTB+vmXUWMFS
1WoY0zUj27M1G8nbZFbmPKzVUEIBxvsfjBnha/jCDWYtMFDAnKePv4sYU3Uv5Rtn
tY2+oNBrYEq1tHkd5pCySUl7cH3cF0q1P8ncBTTUDFu9mo/qA2kNsDTtGmEWwtyC
0tcVMTBJ/OV7U4Czodm7LExH13p+/uSz5Rs1gB5n7L1fFOMQMJYbxZIrk/rhWZHJ
Y/r8TIuk0/d9ASj/qXmXPvEBGuhA9vhMuBlroZ53EGVfBZoY5J+89N7KlKjy5UBe
HbNnYC7AOPMnX2oSucUjy1Z2MUl8gzPN3ewUWoDHUIo76+aES/ywtKxtmn2BSKub
ikkc0mduTyovuXvyRxsOmI2/tpBUTug4ON5lYbfwE8bTVf0keSAa18YSXbNZyrk/
EvyVWYOci8xBUWBbjJg2uxsVrL9ferH6ouNkv9+EV0luzOUauADIku0aKENBdnOK
Q0G48RV7ubZYSzijlsJ/Yfa6U20fbbbhAIVyBXACu/6m5OXx3AhZBRu/UdIDXU2e
sB11IS7q2kzDDguvYFuXf36vg8ZuaOYjlhQ/4UdtBJwZOwO/isJcExzAn4twQ0Qw
0O45KN+GC9xvgn8VBdD1AuZJo3pwKKuPG43F9SZP9Pnb4IeU8mLcv5/lGt8qmCMY
gTp9Zp04S9t+b3p7RdBlluL86JxX7t5xGRXJAgwDYkgGlbPgB+lSdC7wpAmxtPq6
ehsDkL5yOUsCJf1op4gLH5ESK9vuHyYmfxAe63/heaDAdCRxWLI6C8qmhzu52lXv
kAxc8vd3jD7eDw/qe4Ax9pGleJbxc7cz2RoIXyND4qB68zmjbxvFtpWklUyM7abk
/qiO7Kbih/db7j93tql8oMqV9XR1y3K2IoP44m2GlFMjWHQIv05SSyAs+k9bIBkH
JW59/xRiDMUfPdEXaxcvU6P/+md7j0Th3zYkbWJtx5H23JOZg2G7M39mA0aenzUA
3aKBcIpzLsx/DSioOXaTMIcf9KjBMfTRlAHZro87HanFliYXT+23tsUlk6uPwPF3
0imZO74WBejBhHSUlqm+pbPAW1gaktusOlfXwBuEAjhIqAXKatgiMJNqZ1SZurIe
sVtYqeZR3toKtsij9+fPCTGRJIlDphTVbT8IS3Ne98oOjPiKsEUPc1EmWNOKkqiA
sZ0qu8/1xxOToon8Rq/8ZeXAPf9LCcagR+7DGax5iR40c3AM4Ax9ftz1FO+MStMp
G8AuQAt9TI+uhyRywkxU3s7F4H3g5kF93FlrnIXmU+22pQq/2QmagUWEXy4anB0J
GppbOfSZqAia7kT4slY2zso3/qwZRpja3RNGD/g9/1tfHp1eVj3qyDF8bLla6nHA
HrPy0vSHH7cdTxen11HzLFdhArjw9Q8BeQSeV536NTwP3ivC6+7e/se4tvchCSpK
+Oa8hQBIVLXpA4aDzsccXNDhddiJQpJ+v4ciXVMnFQNlzD5jlOsm8Wj/lSxEPQWh
LzMjtvCTjVad0eTAoR/7KJikb4EJwuu02M6voYvQxjnyzlafxLXbvswJY/w7AYDo
fjlmnHwFYPeGDNKtsOvI+aW4z7Pm32WE4w+4Eis6QM9XBSsXe+/M2UrlRFhOHY4E
Lh17JSucnv8F4gGgGYkZ00mmqHcdVY6lc5EXo35yTGgOZ+mWJMVrLMkokxpeuD8b
Ou64HO8vYyu97wHTK6CYRN6D/dV6QP1GFXEFPTjmoQyjWZu+sZWxiN3xs85K4ZP6
5nbgNLznl4VqkTWXSxHsTafawi3TgiNe5HUvpo5/U3NPJCER+YDO6jKEI8ECax7H
Jg9EnA5cOCMF93CL4WpeeT3NloRzf7Vl2+lzeDwvpkeVSbaz34PofJPXt5S0470Q
MDp7IvkgUX7zpNTTKxV5qqFmz/ZfeWuwu0KDjoXk+9e5h/yT7eAfPjhZ3Kne4ak7
sHvSLxS//gTrgzYQLUViJEQBgZqUqkeQ4QzMvkn+Fce1qBgjwHClqiqLnPFF13Sh
IWn5gpyN8kUwjBqCW9vFI95Rnx2ESYIFibbOPtRzZLl/WMX4NS4UKzdGVUER2nqX
YDC2SoaVy6S9maCNpKM33rNSpI+0Q/VzTAoLmLRjx0sELpCNLNVLGOBqIbl0UsKT
AOh1sd6arGWDifYuGk69OZSgqHOMbkPEfdSDCexSuXkGKdvO+/D2Hit9SmJ5RaW0
3QQEx46BAnTEI17W0zB+9tNn/jzT2z3KdxVdTGvZ1CtugzWaBjkhk9tI2OQlAkIT
GMTLGJ7unMd6rnT2ZgHwXTPoXuIEzJt9cwAvBBXKm9uQjnJ3nymq62flQCiLfLnr
7McSuZQgMhgRsEdkYhq4DRl3Ox1rbZ/p5b0k+FG5lDDr0DDg6W9miBV4lqQErxBH
FTtmV0VFZXRLZe3Gt0QCAzAa3wr6LRtfMtPy4xg9KHANMagmzufapDGciiI/wm2O
ngdY6cWK6CKUOVsJH6Yw/f+2EJMg+FFJiN0i7A7CTJoan/AnZt0N3lU6E2t9yMWI
Ln2xFuVFElZ1Go20gsrIZ93QRj8clGbL9V2kxlYcwkw0AeiRwtD8obSeX9a388AA
5UpH+2seCRaZ5tOvf+X7PGVueBv4Tx803oWCNZZSM2sAfGfygkswCIFZrIsCpwi0
sECRuEscMxD1mLFeQQpgYbNekKdZoWdCU+EH3kYLzsBqNPn2AzlbEOyAvSGRdoYP
xiDlkQf7uX3NFrNKmANMZyAygJ6OBvRLWONNfqRxLHygko8R2nADxiX3x6eORsvV
iDb6/zfhuVmJkYyh57yHTvZ4SH3+6zA+HTGPPdo6vPUlyn3hvq5bvifhPistpF4K
KiWb9/5Y0YgeU8bPId1qs5n9j9qfmMVjyRTM1cPBoVsT7TWBtvpcs4BdjK2U2IU9
4CToFq/HS4mOZ7nUCWdXjKF2LiCoEID6r91Vr967VYMj6SOyrVW3iTgv3euXtTVX
rks9cCrIDfWR0WfYrO3fBHFCIThbwFb4qv0ISTRpDTX1+F1ohDo2i7GOyCrGQ/w0
/cqqtgYmH36+GtdQq3pKtUwn/0inSf8EjZxd2CqQ4oExAwVmYi2UwR9KLMZX5LUG
StXZ7I3lx4LIxm/YbmeQxq2TLuA3Qr5Q2YDhKA9BjuCdccNjrR+4bjzFI1J8fCdH
gvz/UHr6Jxiz+Q35w1+M1tr0o2BdKuH0Tu2gYq87/mfi+/gUEmlRU3XhePF5R5Dl
NdaH0ZD8SGZhI+9t/qbEALuROPKx6huAEE+BEqAJ8SWuFvhqatM2ahRNdJ+qcyyt
JXUUhcr4BrlEi7/4dlQ7R5+MpcR+OgZFOJowZiy7TAA4I+bbHym+leFvYw8i7omz
kAiKPsA9RY/cYAUFzwkSx64ItDd9gvWQuwPqqg3+cZqvOi9LRnSHO+nJQ7Th6hJw
d6ETvexqNdTP3hofzRXMu61ArlYT4B1W/CC67nnch5Lhfopy2alJCC9ztrLsntb3
SLLDfCGDDug9842lRYkoS95EAfKB5dtSufbSIwVTBiguhRI4eBQNekuGeOiZX0sm
dtmKPBiQhAmPg9zJSjzcMImEmhly0bBd8mjcutiO9CZFld51YqHTJoOi+7Xohvux
512jG8wEAHm/a7PSNjxMUszsX5HrynBCfNleXio9qKCm1MTs86mmEBy2JldWXxp8
yHOUC5bCSB5P1jRhzCiafT98rA+/PtyO6yU0Tui1/hv3G4v7yyj0xfqj7izQpXWI
NMdGQjvBMeXLqpk04qUkkdyOUbN6+MITL0BsC/7B4bUdHR1vV9nl5Nmy70I3BqVN
qDbtpX5tfXLhoGulDrLctFFqH6p/NhTO2qCDsQ4cCrS2bioCZICb8AnZEj2Bhlub
JbKivlWqP1/LF6X0ErgOJT2TZIJkM8xp1zifYMmXHpQkXc8w1GVIcNjQIOJvfDQf
WUwFhFFfler5dbjTXb8jtLKcj3SXXqk5kdZEQFMtTPUYtRLTesnQSKm2/fGDgIPy
A7ECOLa39s1A1Wk2wJ4g6Z6ZjnRcLv2RWKxEIzMq3Dzc/zu/Banm1Rv98f4pMnLo
3yYYnaupV+geSUMQ2U3EU8tJ+j0v6+uVUOaMFyFgA2Veixsj4xOenl6xhvHwJ+pr
FzKV1jLWr8VhCRXPSkCFsSw9GbcG1Y9X7G15JgMHHjvqfEB87RiPVghBkZIlUj/v
pZlNLWuNC22cfDSfBeH5EVEzPMeJCKprt/mPRV1N3M3NH/eRdV86Bp/C5crJkABe
6dmSNCJF2t5ReqpgTzOtVqG8UxC1jKqLJDIbkvw9g/A3ZAkd3KqKOqe+P3vLnMIH
uYzbN/H8n7rhSdTIOelASgeA1TdlbONjPkSn+9Wq+9MNybD5AC3jGVFoYXLVN+ut
ebyoFl5VWbmGz8phQnNcXPBk1HHGFha2FEbCo8cnc+gF1fict0Acp2AK1xEZ3z+E
nHYHuoGBtaS0+MtfntcfvStncJqC+ec1JFYEY1tPKRR5JEOzXes8ooGXRRbLXRN5
4cFBgLegM5w9syNYMUUPAmuK7zKqIWXud+sDU0GNWQV736Eaqhox/Refqza5Sb2g
ur41xt+z08RxXNRH4+wfDlV/oyK+l4K9R2hJZCSDm42pHTDp38MEgap+ZlxKCKRu
V0Rdp4mSRjgkku9/wgZGMFL0cBo5h6S4z1T6j22ukj6hgw+2yHHvc6beCzI9mRtE
k288qXX7e4uOPzc4YqOsyZgV009TjUIPFyVuZ9vRkrSpb9irzCIIYlrT0jhObJ+A
RQWWpeezkut0EFwkZGMiE6zKeQSj5RTeQTOGaTZoAA/6yux5v3eHreo7xO+EaO6h
c425mNVpfOBERfyG/5XJ8nMwE0+WLVJS2sDJyPSGi3gS08sa6qhb6bSreaWq7KoD
GPxajq9mekVBfeO4RDfyxKBuR3h9RhOsURBvCBv/PUTRwvrzK/LZ6S2G5ioUdBN+
mbF7Lk4bvcmHKZh6FL0NjYrqhM409+p+AG0VcEox2adCjQbHecePnBJlUqSeeU4g
OeyxJWSAzjGi9Njm7OmxkmjlncqY8I1oLTo5P5flgybQAsNNfvPd2mUQGV7Czvkt
CZ1yZdryENlh3dfxwTCx8hXGQIiIV2835bJ10ieXQdzd1oK/24pBCp4tmYfEbxAn
h664jgEQtRcNLCYmItx07An6XX6KQ5UBditaEpEVIcfTPJjXPPxb9UuGyTkZo7Tf
YAYwtqXZ8PsSO82oEYvz/Rtjt4udm7x8o36zgvFIsCAnlEN4k13DQsRN5MNA24/d
Vhu4csoMeX2YRrqA9UHRiq1qrOc8Lw/sc1GUl7Bh+yDt/90DrTgiZaA+sbNIoWSc
uTfJWzpQQVKRqHBFZaR0ZO4aAcSAaomZArvUIteR+TISR4Btys6nklu3YSzRhH/O
yEeturVYNKHNg+U5AQRqfRXMUmXF+VvdSJw0g4VC4iDdILKjS89NZFCSAc1L6Crk
46q/tYV8IcPoog4q6ha6nnri0/kw44jquWiXDL50F2STCFWEIEzfxOnK96fhTTIQ
QGhogVzHYKkE8E8WZp5hmvKEkuqzp0M0e9QgizGpXEzHLIO0Y2wI7AhOeJAicOwp
6Gt5cBiyX3J2he2haQ2uErIREnQU5x1n2Da3mxWgO7y41SWUXYjsHIvt1fIedGqh
5gkpD+cG3dGi9ehBoLmnE0sy9cul+RseCHvtnXgmEt5Jyc0a84ZxUOBNzwQpL0Aw
r77bjFoXSQQ4YVWDZFmYt6FFMoF1nOnZjUdEIrPtxq1ojzNRAKBUELzpQcSfjfPN
L4LT8sFQGGxdLHrwHV2MxKIReeV2lgjudjhlgXRtN4VDTL9HnVRzX3i0EjhORFzh
ii0nrT+nR8aqVhQUjQaKM74CzSd7+gWwmPcjWQ3QTRXLn/FK9NEJrzHGMVVEdLkK
yfZAbpFT/1hWP4MPvn7fnkPV0EBFOAYGdQfYqEY+GHQ3QN4LqZYg0bukXfumh1h3
Zu5/eG8QoSoj3w6Q5XoSsyr4KoOf4dM4OiUOtXTXDCyIfpoIVfFBNCJsUQficXv6
Yc+GMj0/MVUMXYIICnFM5zaARs7nVA85fgEb2tY8Tthsoor4ndOoVlqdsCN50USQ
EKur31E8clans+/9gFT06j8H3Kz5sY64peLcb7ZNDNpNXZ4g/vuEh+N3dEsjakbV
ft0S4ayii8RYXnN/HyA/12xGNIYfCBBCaR4jJ1exh3d/dfU9qPfeyrUnaTqp1Ky6
QIk6lOtiidVcTRNPT6+HbntT8Ne65gJtY+D3YLMUC19fwat1zIVHmZJJcv5IjPKd
egK/lwkD44UxcYaXk7sxQFmeh23DPR+jgdiBFAZQ4KPhkd04PwrGug+biAR44EgB
H6HI2gTrI15XoUDA2uZmvr+JS+sSe8QlkM5I6fl4rtkeSX/1jlv1+qKXQvLZthoa
R8fwVF/hLFu76EZ5GZM59mwSdKV77vLZ/zcWC0CyzCxzrfEmIwkDPdff1CQXWkw5
EhIfzQPtlHFq4vHmfKWCvsEKjcVa3XvT9DzHZGJi4CXbVLnSgB4Sor/XLQ/hyUSJ
1Qo21v6vjVnpyYL4gQj2AIKEkoaOidG5x+QR6+R+3ITVdkaKg7Pc/8x4iR0U74iQ
zNrvveRZ5soj6mTzYPZrQhWZOuQDOu9RnF8phIdltt9JK7G7bmouTExXNjLse89t
5wIcOfcrbT2FZbZCxATF66pOH0r9gLUXw02VlLx6sxT/s8zxmXsO3Tti8HE6QX1o
YleKkG0cRO58uMfCiIBxelg5QfNumpEQHcTP8U2blpf5c6ZwY5lt0kge2vbvd2QQ
yEMe11cVaRUxILntAxDJGc5IXQ3LnCj6QIBOQ9tcAPbIeNaKh8oK7kBvbLaxMQe7
tHOhOvAo+KkFVxgkLgpBmNIcQV6DLf5MPLPEP0gnS8/qzI58r4bk0prhR5NEQRqm
u2dx38owDB0F/K7WKepoS4gXuaKj7MOfT2XTwqi5kBYzB5JERJZqjs6SBbALVj41
YL3k1rLzs2lDaw5YwxaHiyVVqzVvUubUJ+N3SrlLK+N5FKYkiHWQ8D6QFc8g4g3Z
DIJnO6m/s9/hU5xisJkhSWJ9c/zIobUX2f/Z1gRSoCEU8scwc1RbO2ctoKtuZia7
zBpqRzQZepN57EXomIMKIvg4r+4FIESRDPqXeXwPKXsMpkvQah3Z/34aDaVRYINr
QEVBAA+8qMpe1pBI7bQT8Plj3KrVbFEheofIanS+1BA6gOsN+9gt3K4XNSL/poiN
9Jll2PHw4c/gHzRAyO/+IK01/m/KrXfNKMV8KzVcivtfrNbTgpCUfcmD7M+kl3JS
BPVeIVvFhwozLqSrCtp98diFQxpfBifcV9tprdi/P9aCS1tlI6WWx55cnEof4Xtb
fotK4t+6AWT7hb4/fyrpTYQ6dmAGntnfjnCqzVPooHa8iC7URHz54AZT+iGouwTz
YTGu3gbe69iTFNR0QAMyeMKpy5vafjfb3omYgHfSwryymvkmKW9LkQ7/+CALyvsy
VD9b9/7zpq6t2/lihszaSdwGVCSnfRDPRALqyriq9B1hUMc6pJ6fNDI0z1XlAO9t
QN0gl+bFC1uX2RbFdybERx70oMrltg2r4epy2WdZxe7bKost59nQEFPl8TEYOGCs
8M/4jOrGMq4eQ/+QzVDjFdcZfymQaIRSUnsb9KxMdGV47t3e2WvIhWoAGyZxgSM3
9MJxCXaYLFNe5FkH/kBe92H/gXqy76oAp+4/pknrpMf4GEFp+4mUXkkwPnjgrIRU
LMvgrCTlzj1n1NiJtKAIxNzIV6GvUcwtYH1GrRN8Pft4eyVVRNrcieb+DMOQT+K/
88awPFwTA8g890TOaxrTyd2DlLQlsHufqV8/jrhzcErop6oM/+pFhWFlACmF4RY5
gO9lViu6E14JtXW9u4UZyZKjxA58G85yes2K7YKnTmV+KAFPo7/BrbEwrG0IHcQR
QWN0CQN7W1WJGKtHBHe4tjJ5blxCJvgLPOr2DIN0HntAw+pK4tp03bgGSZPS84Vb
6gpwqUZoXvnsyFR9hqNrK+MrNQDiLmT4Rh85BTVF3TyLlSIDOnE2n0DjDmif169V
FGMp/NuhkycjzIhHSmOea11TeColiLoUoUpDwAMyK4d8IQ8lDQMgcXOolhgVii7Z
Owq5gFE5eAq7IjvywwMG8u/N06UTLfFfQKUDO+jka82dPHo6lM1A8UAVYDbwDg9k
Kvz92EBYtAjCt3Cq1eXpKWN4hd6mudEHB3TBEvv8sSs2wMCTNHwEAWfxTBNg6cGi
PMi4C8ldsnsCNgkmw/FdoREVYcs3usYCclM9200qoYxNWemr4JiNWSXWXEVvoB0I
dobClmLJZ3LmqIrwTM5KM+mdAr0a1M9dhp8L6Lm0rmhz5Fb2y2Qp7wc4B/e4IOJ7
GPwwRRKvAhbvOFEEpj6lKoplaUB6JqB0JXDRF41d9cOo5Ki2j43bi8ToaOF4FANx
aBFo+bTyHHX4CbCvuplW2R4JB8lQ+WClzEmWFkqECi8dtPgoX29zA8NQ6bBveE6u
lO3aPGSmwanxQcVzOyOqnkE7mG0xtEsEjWigBjzG39Bp6Z4cWQnaC6hfPWigI+Tr
RGFQLv5G5kBoJG8p+8EKE+gh1YBG+nydq51DbZIwxFfwi3/OXY0PRfEslKjx1/HP
jbnNiTZvUivwyONUo54eIeglQ0pDaYDyuDcrdnG7uN9gDMtS5XuwMONDu0X4oKgu
0AmUjIFcD2TSCy41N8op4EPXbiAOpOKWOu7ek4MSuRXwdiDxDq2PiYp4v53eP2ej
INLtiPGPtXV0Vobj3a3pS2cI8LbrZJQB8RwwPp/W5FdruqgRXyj0ginV5mY2JOpw
O0U+nWovzuBvAPVboEx3mvAggoVzsWzxFErkJ1yaU2BVcHVhj/t1smBg4io7e+w1
Z+8lGAduWRSs9h477bo9wZceYisb58+896tsJoyCsuXQCm/S8TTCkD6emcYy3v46
3LbJRXt/OQFnh2sRXNXQ0EkJz0c4EoPP7gQEUizQ6y+qTtyPrwbpZ84X4xI+E+OA
gipjjjTAriAbhR4I13o3Vm+7paM1KXBTTzPDuptUhHWzPwJer8A1X8DkbKGpThAY
8N0XtkItlZP12SMIMBS4mDgWFy9skfGSjNtsoDt390kjgv4rfGzDb2dhAfzsVluo
+DeYda2hBoOfmt9nebvwCY4xUHIK2gu9CP+bNzYUiCpVvONLfnfWyqiIsDjXNlHO
ixn322Y2yKEs9aazRhVsG/yfaLmk7b4NvypXwNIeSIlLjPvGtbieVIBmqlzdkCRI
2Y4ECgdYCPNME8dGsQanC4u0eoBKdmD5WgueP8xrAf5c0pU3Uc0R+uFZRSgTDl0U
nBTcOqdj5Kz1yrCTyn9urLiMuXKoAMg/AoN5hb8RxNL8kMtLGKahrQr4h0+PUkmU
4mLVCutthTzrXEi7hpCThAZWXOYnRNFQe0ogJBIpH73MgbB7onKTehmZsrVq3i4m
zaNcV20rhW3DL38XYU7eRad2Kz5hnS6GtzmvU+JDVfepjEfkguI2lxzXm2Askcgc
37Nsogo/SLul2bh0ERZwwjVLYCvAQ74j+aRtxF1CbXhtnO9XWv8Mb+dDhfH8r92O
V2ruhPpnfZoaMUxZDNrKM9/JIg9tQuG5SR0WboV6Q3MnAvEZ99+cUcog0LlRnxBZ
/HPhAPuj9pA5YVIAF74JESwfnXxUDEOYN3ZWOn8C7ayUO020LqS5/H4C1yDj/SOn
5NdUxKnV6nWScC2Ma6+vMki9N8DPYbsXYuecHOS2C0PpksZw93VSHr11IlMvBwvV
MfveSvEduNA2vZz/CslOSkGZovDMn52hhj00HPJW+LUqLv1HHoJsAxiibESNF0H6
bc26iFeyoLZDBFU41rNPxXCo7uRX8+GRVEnqMkTXEC+eMb7gc1Q9Y1KYuN7+e+lA
F/YD9DIflSzvRoVXBWgn33ajiwiS8rFzt/LwdGTOF6W7K6/LTpzapf9EyMrtGuNL
z4H2GWRdOBj7IA62EXUqFnjOiZHmp+7BtqxQ8GSzwEDPGxOOhrbetqIyIBzWn7ZO
EEhRgP0Oqlw8YONwwDLYlZHou68Ps4oGV267TR4QhV5gIlAHGp0ROsmYW1m5cIt6
esuSpVPDpOXw5FNmxRqZvorcHiLY8WGKGB8BuDFMeGQLnVssUpXY9k2leseWBxGe
i5wdakV3ucLgW/zP5OS1WGETYAz2lVh0eX0xj3K6bVBFLS7vEd/738X04WG3/tMn
PIGBJClpP4RyXk8nBbp79+H1MYElpGr1SBK693AC0SZJ0uk50R3mGxtmpHmJo5Z/
oYZH0RxSbEIe2S+Npr8ZklvnFviFfGNE3wD/UN9GpYBZNqFU4WEUvJb4JWP3QINb
s31DxpVqKjeLUYF7pdSJuiHFa+iidNbFzoWRS8c2lxwpHJ2D14U+q6R8YkB5ew92
JOmLWUIpHxmIpi52b1UKJ3AwdLpK9kert3BHlC4mdixAljzz6ghAHaQgXTPUIeOC
4FSYiQAH76oNDBxGfMI7kE/+b++qOVj8unO9RD2Wwxd6CWC19U8BnElDZMwxmkBh
27mOKn+/Dxz2gkEaX8yi7XR2i2vNZZkcJVY7VTkVQVKJ8KTXLPtRE+OgE2DGcyPh
/r9w9Q0/CxndX/7qNkkKPjqWQDy6CHBLgC5aUkDpsCVEg8DyMVRMlPxMKzIDCPC5
D3DFz/f2ejCWhvscT6TL4IqySfI/HVeXIk82Tn0+V4uNDvm/ki+Lt8WE2vccyiPI
wDbafYvQsgK88Nai6LkKCoqnOpvE1PWzM8DL4c5k2UvZCzH/YiOMKPpIhaaiRX7p
Zmi6/j+fa3PUc2Zc/mbfijL2ayWoaB8sXL0XIJEZqMpUZnTeFlfbF0KQI2dg5VG4
yCcdbOwW2JrtqyTHFE/bXRiQ6AWkbFH24wWoopgaQhsC/OHjBNji/QjJVYWp1acn
x6FlUAy73bv5kVUkFxqZWzhSsxKb+8ScOMccObhM8PwlAS3lJgwRFwMe0WNRXS11
XidlfLRD4j2qsI3MgkJu1ieVP5O3Am4+mpH3AFC+HgwjloA/0MG1RujXxmpsHMpD
GcF5HxwL4x1qOAF5daNB8WFFkoHHdKEiCYMwvOZMBYMrWy/ULvJi6Hu+B5UTIEjl
TFluqlvFHdY8D11XetnJJklThQckar2wNoWWH8Rw4E9/h33O6gocPmoVaBxtNW0F
t9oCBFNIaxVjP0jo73tw6W7ktPV8yLOKWK98G+gvpkmFw/LYaTPAQluRy4EWikQU
zEn4N3xFKgOk+lEoXbfnzkIeHRW1M79kVJOOt8K9zizST2slSg5VA9xVk4Q6d0BA
vM/LTNuPu1zhiqaWNUXn3linXgCXY+rrWPiSs1k85PpQH71aHwHQRo6nT4D6FjNc
oXzS7U3UL+6dmYUJHe6IE0HP2jLVHqzM8pOhZgenDnJVziYH7q1bkLs7zfB1J/oL
tLJIlC82N/z4KqwGdG36dg9660KQGHcB2lCtg1QP8DiWBA3bscDD8zRUB7PIwbf4
MnCZs2/rOcYsYaWwGLGCrYLG4gRRhLt30W0m59JglhO0OK/IaFNLwFN9rmediYeu
4nFQoSlnq72Ezz84RoSdmKcxmj4HJRAZ2X2p9HfqWCfsbtI+miGKu+z0VX9QBQPO
8IHdcPss9WhLZvvbut3REeO4yY1L3FT6MgP5OMR0gDdVxdM3pwOlm3tn8lAcLNgH
YLZ/ZujrnJA43M89wQniF3ydJueUaHkov7JvXvAjG43Rkp0Sw48s2OiznKEWE406
AbRKmP8DFUL/O9Tb8f3A3GOD0cbr3vo2HP4Cbp/5pK4NXI6Hn5v5i0GqImtuPcbh
nNcyzzSiqWzZ8wliVuZe98n/Q7InPm0Kspcb3Fx0/mwG2d7tx+XPPPEN5EihRCss
4DfWZa76dnH9jtAkspTg7CnpBFEDh3IQwdWE+EgKtdABdKUirG5rez1HNn75ggX5
vADIPvOFZx6gzYLaH3sglji/gwXO1SzcMrnQtWs4ldkYL36WLRBEwVWFuflwsboJ
WLv7462y8W8NSlRvFAG0erz1AaiaOWEcxMw8mfQyUAhidOIO9zAS1E3h7IGhfQ+F
53WMwFUZoM0QwOwhw90zoA8Agy+0qQrjNH6u6BSrGs4vOOYSO9uJtLmhpt72z+Le
Uc9mWx4r3apKDF73gg4AjTv8u1I5jWmWoAAWqSAzhqyBvrS9v/Ez4mEzKw2S1Wen
O/Ro4PUc7RlhUIS1OfHL+lvNmdp+aJudsL3PwBbA6fC1thHMrMl0+DuNlSir4cpE
UN4eitJ4u+YV0A9xS3lbTCPKZQfK+vshsHq9M+4MiigNO6Mf0JgaW6Qv/J5xpl7f
RNRHRd9/qPzLRmCJKHuTt0kMKcWjArB0m4qKVpRTNKWYtwiKvcEA2GoRUqe2/SId
ZemaS7bW8IZ4mBqEIDju53sWKDYBYyl5aapuuGk3bL2PNsAaLCHF6y5IY7DA1Nyl
B1l8bi6SI0TBSrStvk0zZOcQLzZ5wcU1/d+gMN3QjlyGNQzvU5OLSOfZ8t6sLYUP
nlhnp8o+0ZtZaKXEXZQkJ6wFisEEr3ML86+KdgLvMbPPkxDAvypSHAtAWDok/gGh
R2d2Nlby6ztQzaB3rFGTjevV51MGcYLv1Wibaw26FQBDCPDFovNXZmerVmP8/11+
103WYaDh3ezW+4XFYgvTB+Gy8oin5GY1LIAMLffUrX5kEkcqq8W1klvSlhxQAQLI
/DhAf45oxR4v4HA9hqwfiGP3ONziUvL8Xc6/dgHBGRlbn1ALX7sheTNohF/gb2Qw
hPN+EeHMrSgBpnn8XLOmoD39VjiGVd87YsrLijmDIZBF0hVWke+bnahAUYPKUBin
HstY8OlIFRbZJfopNDV4Nxh+p22ZB60r1OoBFxBdKKqOmzBICNM3b17DN/Lh3JW/
QYTgQG0cFJbtQ5gIz0b05gfWadJOKUCOxfE4En3KLnsNU+AHit36oohvjGB1IBu0
z7OaNgdih8qDPjViwm6e6s2hkAP8eRiiKpUGMPTcOFwuCRjXC1x0Sleb4NxljW8J
H/xY/4LrT/ygky20Rt0cn0S+k6P8KiHmQptFKKu3LbLncTIR19DvOrIdsoy5S4Wd
ffO9tNdbcmptc1EvUIMlDvLpiipivIjQHH+6GkUH1BFmPe/mwZCyZosUiKgXXKEf
mnnFTjHyoTo6Kz693AIgytCYyLX8xwFy5GptVSKoWIwDNL96psrAPKEQF7dK7/lZ
JQ3SWToF4fB/SY56TkJigaatbOdbvK9C+8N8bAMEfrrPilWjI3yHqPcmlmmHvnOB
mowWmh8FKQKismmu7fnrqy8jCy21qmLL0qlBWrugtrWYk/5LmQ7MR+GEhYlXDrO5
R2Ep+40Zl0gH8V9wGUefd/zze8YKK7UCZyRTgyKxDnBqklMM/xzqN7dMYnzo3bMR
fXS5piD+J9Tlado81spXb8t1zo75bDdzK+jEOoRmnx5S1dDMX6AkNz2uuMmugbp5
il6ySi5GICA1lrySY6o8SvERiMf00i+LntmTabtpfvhyht0vWTbs0FEIXlR9to4O
2nMbJ2b0dfWEMABMq0GSuUrT52pFCsyWwW2fzHw7vjm1lj9bFXYPMrSV+aUMsmvU
j58ZGIFmp9/1CdhhhD/oXkrijYexY2RJuX2vgFwWMUyYY3i6azS11yL9Rq1iuQlI
JYZWfkz6qrHvfWMM1OGqjffmc4eqvLMP6YDzO9QH91es06iWGeeSWR6jVZHmxuow
jzLKbMl/gGZAibhrWCiSPCMLKUUBgACs9eSvs9cPpJKAhPR2DzIxODhO3gVk7WPP
qkLOUUkJcyZgY7HSe/7pZvHBV84XyyFDy4RJu4cgBHoZy5PclQf74GyIYbcZRdZU
qTY11Or0HMDZIkurg9QbOvp3hV2Tyg0fxqVZ9YPQT/jfWktF5IuKVWo4Ku3BxJ+P
n6+RCosJAezfxH+X3St1vr4CgS+jNmZmhANV6oJCw0276Vt4oJ6epCof4rQZM/Us
A2fzjDqZr/A8mbsl9ApwJAL6Pel83Al0+biXYaQHPXwtfHGpzM7xDL6Kqfh3mthk
2Lk+9ZsEmFYoYTV19ESgccWr+Y212wthIzYxBH/b1qHvN/98qGUqzOglTblUrL9I
XeKXM7qUi+dROjCqFPyV9csRL0lZWCeR9yFLlRI7vU74ipYx7/ZcLGNw4F6VReIV
IAz0m3IOKR0tlfSnXKlI8qg2fI62nbbmFe4DOyWlfzzbGtmXmp9KydEHvOuHgwRQ
ApypTRANW/AhW9VsTcslXzZd38wT2A8iv/qlpYEZScOxUAXJBpJGD0dYROmJ5cG5
TDPKQza9CyvZgNG7oKJ/SqNtn3U5ycsseB74SHX9vlS+nBRnKZfjm2G4X+UwYBPo
2BI/ZlgsEC09seJ+2EUECbXDibL60D8XAOqhCahZ0UKLkhRvHGFd2dUekYQQq/tC
LfLMFTdBgS73d9VgeS5Taof491h830stu6cb2JOEQKFnmemS1VO8bqSUdXY1SOex
IbZplZSUFtbctM6uTQerwCUF3peX1OOl0eRBz7X+Gv7JUf2RZfQSlNurRtJUQqpd
RAp+w1gin2vWLbDMgScuytCnx+CHcvmDdQ2gRi7j2W52RQuj1ZLiDGzFqJ1gHm6C
xjjfnnfWkY4M8/on6n6bgVMH9EgbFW5xjzmbTRW4l0mTML8JsrI71s+XOwD7+d7f
DkV0u88gOc6l9u0gB8RwpaxvbMY/ANgoeNcKhMwm4S5Ntf2pX4HmoesZs2YRP0WE
wJCbyogbBb4MKZ7jBQROV5wjcqqXFUbKOsMa8TmS/rZz4QnpVanS/IJ7ogq3BRRl
4xZJLC18M7pbAy6XdaLoaVH6+++Vbi0Tnx0Cth7IyUkfkfWYh4AAwOz9hw4hywHw
8P7Fx6NGRoZ/aaFIOm1T61Eo3ucVL+lS0rGBvJ2jbjKf/0vv3LAAZztFumpN3mMX
rwHSI8QiqGOHAS/qlVbIvwelxQscC4rR2ofkSzAdS921Jqnvv+Mi/2LybulP1zRs
MsACH6tIn9IxbXwxmyDC+CX/0eXSGzSaMDNMWYuzWh51h0aFFAcxSpKRBSjMTx7+
lK74zBRRko58n1uqLhPNh8YZXrgxjmPEEYmaCYiop7TmfUo0xxAnZuG525t1L5nz
GDIzOYtvymTun+BLgDEqN7SO8qodXaHGiK6/7mjincTV5a9fo07um9HE7PgKvcTT
vA0jXd8AM9A2QHF+YLeIBqr50tGlT2bpjbGfcI46FMqnmgkpsZhmWztnZUDrdm3s
L747R1p09+fX4AKZCMMp2/kKuxvvo3ufqadxMC53fTAr2dnny2c/SeH7UY7TglBL
M+Xx1JhQlkwp2JC4NDjjgh98EvcYskMzNLvGP/UiVzjvfW5/TnT7+gAoNCk60nqO
ryFTiuI+7TQZdmopd+obGJXZeonlY97w0X9t3soI4OGcHk+MHQSsbeo3A99ba7p+
24E/CVRcd9WS6js13sTUvdWvlqIG8gLpxlvzteiqN4lDHv/xQfdfCFs8+G5WoV18
10sc+KynxSwcP6xZ0EwyQc6qscGgrTbgX3EFJ01crD2PjqUCjFeD5IdmkHHkxB0x
EImpXZYKnpEDCPSK83BT/2K9i8KbjEYwRwimduxm1E0+3it1VeFkNYtQX7UBPJt8
7i4zFQ3Za7quRPtnUG/CMfCJnQM4zkQRtplP83A1yytm4vXsM/akxaBWB20j8ly1
8vIc9u7ZAXR93u23ZvjUdmbx6b6Pf6r915hABmYztxDKuPKNotr4z8tk/iF5ZvBD
dJMx3ZGwS46SE1l6EaruuAOW3xCelPxIzGV6/kCzeiZ8IKRI854XJOlKNwqfzNIk
mAinrmX5HCRQw1VxEkEWbJ7SKm1mIVHH0R7DkiF/qhdnMvv/oVKff+qNHWF8i9Ty
lzzwQ+v/+QImaZ7IH8eJSk2kYKzp2I4uEDHZb4nCwqU0wwdeESbqWHKLZZu07xTm
M0j4uUpqJTCoTPNsbKz017Gpf1sSD2ZOhFCd9GoyvoeBO5vosKtpm1+9OavgUjdH
axlXKBNsNgtSu7J8DSj9nzIVuAT5WVgUqzAk1DMqGay04SqAyfXcdE4N7ZGplku7
jEa7dSqcMWun+A4fsnUj8ToLmuxZLeipCLoTqIAgpR7dfLULAyGGG84pDTQvNqB5
1dWX70Wz2MghN280tbk0/IJanvRMy0SRJCbNTVXozBD3sNp5GVRua/lHlD1ic5tu
KKMXxpdoXOQyfiMzdhR7y6tKaq7JMZBqEi5uZCHQKHgwJI1qusV0XBmv8zN/iY1y
FZpeb35IqjaKlOUkdPAj9mvwzK//bAj/cUNHyyXLLQlCrXw3CRRiXAdXsJInUpYp
AgmNUW+Q2N1i4W/x6r3x0EgGy55ol1PggLF+Z26Fw3n/xCtMBGVkFcXId8gU5woh
dieGJH3gehyqpS6dsZ81i4FUjQt5fIrpy5P3HR/vIWJXQj7QkVH0hV9ICvperJ3k
tIJGpBlmyVZguZbfdFiwFv9LzsOoGQ/AStBQ+vD20zKJKETtkzlN3nJoeZd3Xfxp
BG2kF5umVUausftIptIqoZBNc9XEEsK+rU3Q+gobsPN6QloNRleX4WJ2yru80W7K
FzuRnmrFpUyTX3QJ8m6UeHcPWAdXtaoQfisGVxpWvpSMnAm0C0/tSRY/kZcLBYBu
zzFc67UDbUe4mCTlbZuCTmCttFo/knALpXtWkrYhtM/SZMp4S4ixy8FcvzMVwc2a
1B67gNllJXVKhOqg3D+TNWkMq2N/L8Ja/bmzfMt3AdyXBnTgOOjGzdA0JFQ7NKF0
XKof5QD1kTo9qG5EKpXtts0OGL9ZoQz4X2kYind5jHdCMJNGL08t2GMZOvjEWCCI
JZV9h7RWuum3Q1EY3945c1QO3YkuzC5fySg67gH48UDiXiggSIZpRYa1m/oj/PyX
YlsFs1BsW4lIdeBDDDWN9BmXhOpxX+qP7PQ0lRfvSswF7BCp2gignXjtGkbjOiXs
GJCH1JdtEcGwJmD5Z4m30Lzi9zd0bJPD3Z1kA1qqnsgRP74XxUXTFs/o+b9U+561
XC6nhA6l5wKEKGCDlBiOFmLDukM8x04v+3owfnvN3p2tZ4RtiVbHDe/Rr8MRUFwg
oJPw/c5XTEkV1T9PluxsAHsDt5HfdTjvVzm2E3LILCCMYGBlkQrBL4PUA4Lrj9Ec
lTfw46H5wa9qMbckRkh1D7adwV6rQYeGyg1D+KhPPykFBL21oUauy1s4GPij6bvV
xS0TNcDFf5zoNO+UNRiyGHidik8EOqllXlof93NWMuoMDgtbD+p1cJzQUWnbc3Xr
gCEFLoj8mDFXlLgLtOjr3h02xoPjzlCKUrzfe2daaa38pGMddjBUqJwYTkpQ74uJ
OsszqxEPSxjBcFRaU7d7JLcBIxrfDZbMSA0J6V1JgIxHNvb7X8kuSM86oOPj96FC
J5vbzkji5/Ais/bHKl0GU5IwfY3yd5Vm0cokUywhEK2jo0nup8r0E9CtgitSPRij
D/dl2EUXehzf+HxF9PVK+gitnD84xMYU6mMJH2uRw43kOl0pxokNf2mY2764fl4z
LwCtNTPQSXlqzdAPMOnXGUYHcCpjw0a6bkC9IDdAZuHn+RazkfPFSbsrh81lDL8z
cBctTn7+CfSQKjJCCXVOWwDn3E3LVJSsZnzLQ860iI7tyNisMKFG+xagMLIm5F6L
4EQaVvb9oEahkaLIcl0MHFgYFTZxnHkYUO0j5zBbD9e4ELZ3IkXfbfjwEDOWXV0l
w4bdqlg35XuHZf/Wwh6aHmLLXRjl8MBFaXPb7SGzHTxCgWSA/sDvKxpseey9ftPY
XykM+CJjO001MLqhQzdrC9GXY0OEPr3aI4RR/8idd8wc5amk3iPb+kvVqbgE5ZcO
ftdflbRkf/iMSupFXQzYD4LVwLeJsiBm1e5YdrifkYWGDHOEKMxn8qPCWele8eOm
T/vr9OYay8T1WwEXzqmsDoeJcC9gAWZWHHazETEnqtNKBTu1eNZ62953CO0ISR6V
6iKu0S/aaAtXMGej5PDMT6Q86sH5RfRCv0OPj+V9HB49kpI5/PRNuhBDMvF1C0nI
gWTpsBT6EsVzQ90TVeKC9suto1OPPQxfjfOyOC4KxhOD38Oz2kJ1nBMdTP5V6Jly
XOT40LLlD8TGEko69gl9Q/3hEQJnbFuMgR3E8E7QWCtEad2bydvztM3R7othUSgO
+0lM6Ra4FKNaqf3iRwFVCykMdvR9/I+mtpYiBz7gNJCuR68fA4Vu5xBatr1ul66O
R9BOKWioccoXMJ2gBHpaATN1+IVjDNFl/EtTVGTXILgaC/Cw6tDFnstACJKECMqY
NcE/aPIXplZi7JvKd94kTqVc04u5Or3FeYYHVzYRw+qAmz1SLCPV1/wanBrhK6m6
o22/dmNnPrH9HtFSCDA0dtVBTP+37vpfH5OwcklVif2WpBQPtaYujyOTEHdwLney
glCQKyqr0LqSBHYWn5xNa2bU3VtLdil/J1/kGn5PpvqdKBnRlWTntqbP3JUPTiEM
A40Hv93E6OvjCSDi6IelA11WwZUWQbW+Quu+IWMoVT+rvE6osa5LAmtFRJWsGqah
5csOaiWp/4SuvZtv8vJLAg==
//pragma protect end_data_block
//pragma protect digest_block
hizVJWVzUlXXBIraJd2ri+BOgIY=
//pragma protect end_digest_block
//pragma protect end_protected
