//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
AC3daVI981j6f8dKbztGO6WfR8gtGF/Y1+xDxnMkqYU/yyQosJACelkAqoUEU6gY
YCmhskU56Fo6d6KWiX4K+A/SiP1ZR3psLWw1S2wNfHGoZMuEynMwz7KwSKFsKVRv
Q3IEyNMqPO5JfKzP1XvwvPy2W62bKHkq9N+tayOjPpNCp2pq+wwJFA==
//pragma protect end_key_block
//pragma protect digest_block
IM6Kn9xPPQo7idx64/4ugm9T33s=
//pragma protect end_digest_block
//pragma protect data_block
INYa2vynLN9bWy6KgnywZBoQ1zyUuhaOgiA4147erlnIBhyyaekKKwVnUTaBDHPl
anhB1H+HnRYnCuZdNAo63Jn9KdCvu1nZtgUz6aiDAy51/anL/uAYtsYRUkOUsDOG
QryQmzkGfmQ3aVSXYDo4u5QvB949G18WJQAfJmO4TURtqj+mJzs5lB1NmxU+wVo2
Un9+olgLgLXkT0vZdpuDpyffTZiZ8P5w+YLBpaDHVxPyWqg4+YpVmO87P+3qFTA3
113nsDFQ3h5H8hfWdmC3gllGVyAo6kxhmbipc/KjbbvUaxsTR0qLl5rLAwpd8mBc
gqpBuOKQFjZz08VI1I2D4Q==
//pragma protect end_data_block
//pragma protect digest_block
IdtvAGZF1YSjHqqexpX4e+MXElI=
//pragma protect end_digest_block
//pragma protect end_protected
`include "../00_TESTBED/pseudo_DRAM.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
Yte3Duc88M2i9Y6ZS01ZQZbWz7qQ/TpXtLPWJozOofv1m3Vg4yLsuJjpQz8+txRA
Jw9za3YURR6ZDBQq5RRR33bbOC6aUdXjaCKj0jzDXZP0kSEcLgHfpF+G+aQT/E7h
oQNhvY29p8NCXsQ0aaYoCnXFOFvqre7cdTR/ZTXJEdMniM3UCNKmWg==
//pragma protect end_key_block
//pragma protect digest_block
4p+PEPDZquWTRj9Ap3/nEh0KJHU=
//pragma protect end_digest_block
//pragma protect data_block
N5WwoxuBb2d/QExIr55gs2HBDGNPWYOZ9stWlHlAfGAL3S81uHW5eULJHYeynqOx
dHwQRl2S13Uu1Q5u6024jcXtwtcV6WNxoODVAE5CENatpJqVAfxDW7Fb+BdhY3gx
XnxTUjISo9GcXW78PFH65lm+mL3ZKeiPKnIV2L2JrrLjbL0ADg7YKwdZ8/9kkE38
eHlNFtu5GI1wACIbMmaPlxj0ZtAj6FVUEuQdyzcD5XEq7fWZXAjPpSWIyPUkFu3N
i5xmFCsNbzBjDSjrbzBmR3n93h+F+6i7OVNbs/+vWezjHaR3l7Wbo3jOfboPo+rr
Aaq2MlDI8N8HtbkvPRoQ5Q==
//pragma protect end_data_block
//pragma protect digest_block
k01Cka4Pcusl+QKdzip6tcr654s=
//pragma protect end_digest_block
//pragma protect end_protected
`include "Usertype_PKG.sv"
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
ykEAAG5cyEZNLypqh391XK17QoMmLvq0e9hVsccc1dxXUZzawwXqI2TOoM5Mm02r
XMhpIet9EGsf/j0XxbdLeu1wPqhYnDJedIV8prBntASVDWyxmwkNqt3uMvgcGzkl
sDEHvA/aydjOB8lzqWMITO1TV/DAdscmnlHkR8IiJ2i0OIDca8lvoA==
//pragma protect end_key_block
//pragma protect digest_block
SrdcKQTnB3unmY6OOX6owA043h8=
//pragma protect end_digest_block
//pragma protect data_block
Tstm/OMUg4bMHMDL6xaKUI6ifDdPjRJ5RyTYlUgREQXIkUMuY1vUqTzmIN5RfW3J
BuTXOHJhnDKHWbP7z2nrObuuMQ4FMouyLy6Ym+XnTTXQmMFSbkjn0DxmGn6sTUHC
ZCd3d0fg3wW5lbcWR9jXUUU+gpr/bobpq9QwNJ04N2YDa5eD5m0BhAzhKrXkRxNL
SKGeTSdIKpQmu+g3Rwm1MTnCbK968eq2KmH6HEePjCgbrqp7CSuaIPvQ2UwYKFoo
AqhtCILV6JmQdK5mWeGrBqkWtKD7VMxn1r1Psep0MLAMkGeWAhAWpFKC88GqKGb9
uOUlnT2faxqvyhv2SFT+OspYPumAzMaSDAFqBEE9n209ZHCmaD2D/kEMgPyyb+hF
3q0XIRdlcP6XHl51IOjKIUGTVPjntmJu6/poUvW5FRbulHaSDZIxXG0ksw6CoCfS
CXarj7WBqWx1I1uva9oE0cA0hhiORJD3SER9kdke5KD4awZyeGCptFPDdbdpQ5F7
tckQYl7zy9cJvHYnUA3gbssxeLTLzoKc5VBdCzvKuucUB5nqF7bPKP8+5ahzF6OQ
9h4iTzaOLiqCYU6ckllpYYj/vm6Baw15BIoOcBCrR+HlDaCK3SwJCVKa2q+VG+Bk
nDrtTc+JhtS0vvW/nFP0u7oclRaMbL2aBfUcdOdO+RNmxNSf0AUgFiF1RFpzQjes
gnUr5qe2XQy317wrEUFOUDzaJJHruaii7MwXZ9EWqy7E45auLEyWdg/MAITCPIme
EEznLVVw8LCQpOBGqdzNWIzg5SFg8zvnrN6mq1p1+V/8ii0oisXY1RbJgMy8Hqcx
gKOKzML1j0if59SMjivL7I318OlgByam2r7dG82RS95gqtc/XpbM6ogcKX9b/fRx
XcwP/u11oaR9eoYTzxJmLt5VxviM5q8yNdasGWSNUZYj7V+iz77scsNCbhN6GqPr
vev3UpzvaP7az/eLfO+TSPWM1yjZI0//MQWY+Zv+EvAxF6NYfRprJXuy234H8A98
rxfAkG6jeTeSnu3cz8ELTE7YJvBM75U2oe1Y5zjhAit92VWsWCrWS4pCollkzEp8
BaYpUkeOkA6osADhAEJdSTAbAvKzYEfZjXytsZU7XZFss7N+N3XWtfHyeXqKNZ22
1Kc2EcIaVAuSrMa04ujqs99s7fnrgcmgmQreUbVhj4qDU/41/SjR0le8koZQVxlw
cEH0Elcf68JLbf4N4UhFQerJJRzdFxFhKYLd2x4VKXClJ1V3scfc2aNX5WS9oNSs
cMSIUH+kkGvq/2DzHueNhv9LjSk49LSBkDJvAaWNpCFITtGqJoFVEFTwC6cXf1nl
BAfyWQ2+vVxX7eUVLfuvYqKAu7gFKcsIjnYLPOA7zLIyzXZ+LnralAJ4nJklpden
huewWHY66O4Ks1wWIssTFOMtt6Q/QqckN2euEash/QJ7bv6Dxwin3SLJ6gl27xUi
nAF1NH0cIS45N4u1m5bCs+OdE5NV7dNel+tuk8j+jXdCiyiWTAAWNmqMHQx51vf3
kZmgHoU6HxwnjU/GyZJKiopCoN0kPUkZJtndKBRERW68eHloAnhJjTRZOwjq/mG1
EzgFcLEDzSlHzO+uIN+5AuVmCutqx6gDku6eToq6soG0KHQfF3FdAILEyWUovWp9
5nG89P3GPVyoSsEVHNgneydmuD+/gRDfcmLxZgI0K0F95wP8ziS+i/fuMov8TzBQ
x7+OUHxlIxaMrxZHJ73FcVufdgDQPD7znqHxKKkI3W8WVpHgZGB1cZqHxkBf5jTJ
iP5pY6GpFsAZBUE24npw9zxsmzpV/ujCWMM20lg84qULFplZ7ogf5dbulbILBuGy
ePb8mw019afVHe5MdY43xc+qQmCGDdl15uboj4bYECqmc9QykhYGFmNPsTiIwjkp
CklGbQWL4UA9vJZJ4GR1ScxEceowC3hUBs/ccmDPGOrWwYoR5Y+xJLAXt/q0HSRG
Afhwi5cOQEeNMz0IpZk29tRqYxIZ6kWMW5zDt13PWPFDxBukemaRjge59C5r5ofL
oGUICVuhRMyvGi7sq1YaXzsdf/uFqGzzt9cgqMja9LJkIBWDVzF8gsT70uR0b0PC
Fau/6Lnat4VSzbx8JObv6KJ1KqvSgBhEHS7WVDFcLTBuDTneDFQL3TI7TAB1SxXD
xk+T8xzY8amdvIv9xGEU+WThxpEtdchi7BqtWppE6YO4O0Anz9vFHSQQzOO7jtkE
3DWQ0ZPDg0AnuoZGpyqaE7Kz52JWsXDFdRzBOt3cyXMXrEvVs95xGCL3CrFmhYJJ
SBArFctcASs2xFl7iu1RiL/CKbNKYkVk1U0Bn+LgrAN96je8RD5pEK5ThvDd2K16
Z+h17ZSYnDTJ7dTZEZN1p3bFGInRs2NltLYsckePD2ZkSBzD2tkyLZGj56owvsOF
rabYY8I2Jl79SGcIlVVjdXf8wOR4zHVQ6zCU8z/oedPX9qN3q5Vy3I47jP+w+6d3
VgbWsZltTjFM2E3E9+dVaMfUskI7R2naEC1kBqWg0CPrbXzDtG9jta+nZMLjgkHg
BmOoIXe5sP5FuAqQPFpceUGHocl9Q43vGqJSYKFUYj2amxzzsXdKIoU33gncDE4M
he37aSezZGULqF04Szna4nN66dg7IpDdtAp0lFkLo1jKiYDrkf80ZUKPh/mKBT67
74zIZyYbIfrXHSImWNrFRx+/BCyNPUrJ02Pnh0GSj+MyNOjuGA8DRicN7WuyIgzp
PQaOeO7YYJusghp9l4Tu1VdVjVF8B1kL3rAyPFwGaZ59kyoRSkbd/P0L1RDgT17D
OwNSix3tFeNi10dcigsjDdeZtmEiZUVmf3K5JVWctaIfGJQ33ByIB3V1QLBOwRgY
XDGu46Eei/fgUpcIr1ith6P1kK8drbzYTN+JhpLqT+IKGAwj8fns+f/rRuGMJM7F
hlN+vB9GfofUPk2OhHKIw7s2eTGV90+bDP7lLwKz3zOV+1NgbeDkbU/TPSaXAGs2
jcxNaYIYNRFl41kj9bMLUC7KkVlSnxLIWixX/ogM3RnOJDwRo4oOLHXnDiEBxnr4
XZGK9ML5H7DDsDN0yYE7c3bvadwMV1TWpglM25Z7X6UjMOW9x/QEDnObV+gSZ7J0
cQyrIsVgqb8xcj9860Kfgj/6FGa6ZbHPRpFdtL1VozNVLJaUVAzfqDJ28y/kKf68
SD+ru21qFUln82wD5Mwa3vDARPWzZeNpnzwbdW3n8wx/5N+7ew74w/7lE8uHfHgR
Qxs9RqboBdWGkgVYrUsfezKLgERtzeSxHPoWtkIjGr2E2fhC/D6Uw3f/oHBj2IAu
xYoBoY2iBA2EnVQVA0VEfkrxpGjzyyz/5qH8Ji8NZ4AvBfybr67pidbcMVuubp55
2Bmm8D0Co+c3ARdxF/VsJxGSCyyZYC/wGNJ3kEWsTkjv2UOTDyPUHcB0WiSzSnj5
bzaICj2YNARyt+/6xllMjQEBn28gkOo1DFrMz/CmPNE1xbi3hFTFqtMQ+eY1DYVb
VOIG1GiJ8cIQ5PNwbupEtih8XrXh2TN2cNQlPIl+cmDb926xb8ORon3Qv7ME4hnz
ewj4b9rWCUbry1DgNAOSiy0c4A4BwYoKuu+mk+eDuSDJ7U7ldNvnDHXNRDi+nM4I
mKx+UWoYIXzNX52b8dy82eHHDKH9W6ZC9PqsNsnv1ZAF6oIqaZA9hnGEybN0NL24
iRx0FJeJKs5J23xw1Mp9FxyRoiGbvv4Nfi4pNITcY4PbQ6+sRRVNt5bwpgG2KR4i
SGZ47TzTlIw3MADQUBZq0NIapqYvUv67vndraRVF3DzEPUKVS5MjHp5HI8KJSmTt
rMRtP5S7nYkxanjd09oBgaJ7bd16R4XuRmgEHKshF/jIRNi7pqTaHEOma1EhxScW
ddjZdYR9GCk5jozbnaUvP0RwXocUPXdNCq2u8+cMMsmOcTvtGM9N+3bCm64AuJO5
ANzdggLISRJO1Qg3LiDtyHbXSFxikVqlRaP+JFIFqpX1njo6kqKv35mhVXAAYYje
ItIFwsg0LzulubDjfaKst55//x8sZ0Nj9ZZ7NNPrr5QMv/exQLcG1DxVSEGY5UHX
2pnk1KmYq7e6CcYZfGsrhnEXeVRdYfjDOK92QQGAhFUSp8A+rG9cF13e+4S0zPX5
QOeBTbERIn/NGOQPO3hNozCea9U8+Tn9V2RW8Mj04/eHLAcLuyq2pK2Y4zDEC+VQ
59CYY5/zBdzsKcCS0WH4rD/4uortRxhYYjRok+wyiaILdklwWDr4p4sX3DY8q0OZ
EHuEhbczlegOXq7tkTbyh/qU4aznO8UFGXlMJLIbOzsKu6G7YtkCUwbAn1u/+BiY
QoExI8b16SA1L/26jpp21wdHPnuyES4cO8ytlsSNYkIewfbJhr8nBsRcYjcPfdai
MIVRaQTi7X6XTT95JKyI34K44NdVQ+dNvTVDJEYdCnFVhz1MSMyCIDgRfXb3vgeO
ahhfCLV9r00aQLD7vFHwWVo7/Rj6jq+b0T5lSmRZnGAMSyfnb3dyx4bpiNjGIQFW
YV+wgLDZ6wZRqnBq6fqj7Do0tGq6g5Sc9vUxfUte28odDeu10KJaLUprurJYxOpW
AHEzvXILZ7VY+QPLGtuac/QQOyhnie9cMtW9L2B/nDVNGAJRi5C0uzDAAMghuxRl
JM/I+eYXAwXsdLnE6u4r8xjD/Xg2XF9DjQGrmpr6bsPPo81qa/E5yzfuciDzARX/
kEOf/XPiApLW+lgUmjy9nveY2LNhbr24wTEf+BTJL2UobujhOKd0d7ChF+erwn4F
6DeWRE5zDLI97x4itJZe+mTFrss4tcGmeoDGA3k5oEU6y4g4LU/FpdmV4RxGEK9O
72WiL9Lqj8kkSxPtUSfZqq8kqtpku1Z2olnNKLkSd0FubsMlwfnAKvW1dKMVOfEX
hiZXrm5CHkWSD5T769AHGv4dMNHVdLCTrjOvzI4j3P8FfsB/GvVWinmu5lH1bK8y
+5UCpyX7kHdJkNYiI5XUFKcUPYtyQzJ5kwoXgg9zVpJ0MolqMYxPxb3Hm3yVIEIn
S7rmkOAS63g9JMPmhzv+wzQJqo/Q5DCt1PFTeBASdaHxPOExOwmEJTdOm3aOejmN
EMeiY/cwITSdsB2PpMsQYAPz1Dw36aACxytLe2mce1/LxcpniNQXKQkjLTinS0zW
P9itH792QU4knBQIZkLWTON8n0zRldYgWHtWXj3+M9rEMNkUb0HoVMJKDOFKTpOt
eSSrcpQvWDbiNeBla+WRfhjUeFYpd3uWy+uV+V2crQa22bLxeYGwwjBZCYWSmcjw
kdGdg5VpvwE1TZIYIsei6ylr+9xuBPoot3Rifydmqcklnxz2KKhVd0B/xEgtzhxA
eTeveAOVKRyKLenyo61fk3PxdPZgJ/jRnaBZ5kHUd0wuQ83HPMLA0svB5RrLphle
VDXLlsEEi/y+TFXa8OiV229wNXKF6VsxhdmhXmGKLu1Yt/fsT/h4ScI+zq0V0hDI
W2XjwK/Y4bY23enRuCVXHhOTopGYoPPvokIQPa27xLKk+1kv78FPwNQh+omEpom+
AievWd6AOMxE5/fJh0yAoWPn8HhY5aCNgNm7IPctm9NNGiF1JV56ewAJ4/BxtFYy
NXQMNcIsge6MRSs40nj2FxM4KmVGhg7C6Pe0kpXI7EtK7HvltHgwBhFNyqhkTnR9
CgmgIIvBo5XbNdmS3QNgIRMksUmR9n67A97EzKHZrnUQ3EEdfWMko/tvbNXwZvi2
3Oq2Ujv7kL1huvd187mK65vJDfVuYzmPJ/sUtmlVXB9V1GRyCWPOb/V+tPHCvz1B
nijd/QVXNFbgdI0/OTKABTOKu4BxPH91sUgr2OLryBsvHdkiaYb0H4hzyrc/VfVE
zIchptYmBa2xCIVZneDOezP5kEMdx1o7LOYVS7TD5Zoc5CGnz1tHCAE8ySIqkqaV
3lyJL9fewJF/i8mLRRzGwsV6NMHP1J15DksDPEZMHg/ZRaP6h2VR5hGmscc65WyJ
y5LFPCrkIVsFSOoH+Up2BcSmknX5wg1pY/GVI96li68UbQryKKQ95tdfSNuTHBmi
AwpzZtdLL7o4p8TGE7FLhCDMdv0qTlmWk0Pb4LmsDKJwPxxQ9EwfLqBy0rudaTKT
Gf/TPUFJfbum4FKcf6+h3x+LpNnMsRsUpoB+DCn6I0F0IF7JbfmxT93dhrKM0MCN
ia7M+wAO+4iJEjnTqd6eDFuptF4nAZ6w5HMlBnl/7kKl0Yd8BFDO6to7ZRET9CsU
uzNJzkoHqR/XEOe/tFZ9jqAxvUvFunU6HphGYftb00paaWagzL9DGiE1Gi8eU6VQ
I4h1iqsazc7Ptg18aEBOK7BemKdYyepNGksa30iLUa+A4CCkuWmPp1zU4E2GWp+l
O/rYxK63T9tVcov918rBUEg2aJtkRaKWYgDqwI7F8lZHC2ecmi+vEFy3oRHpMfgt
zaxaxnk2mPrYwJRaWiKqeLvHCsfHE1Qp0Q7rCKTPQQ+oYYPsvxBH9ljGFThCAvKV
s4ThNuo6SaVsC5dipLDc8eI1VoqweMtxUjFupOM3WKLju2p9YKhu+pZPuIxYbTZa
b0cVxOp0VTUeLsN0YkYz8FBVCG/0ovlStJWHJP111J8fNclFyScOPBbQHkzHCMP+
xG5n/jXTxZBhx6ePBCgqZUslJiuUi1rvSegKxsLfTNPhiWMIfVqMZk1faKjmlrNq
9I4L/4pSYcYlm0T88HuYcOV6gUqj5s4M7TfCP+PKXV3wSxPbTbOdmZWLF4kWI/wZ
1Vw40ogVHX1GIq67UOm+A/NZAS632QEe2xcg5d9iWFh7pOGzkUD7QGgYYAqfJpvN
qeENjIBeXnaqPef/F4CMiKHicxLdnlNd0ZcuDC7Pfalf/sMlxJ7q9NE/557pgiEu
qYkdd0mhU4rG/Jg6kO9SE/VrlHdDEAlqISE3DR/GkaXep0F3NXPPUUjYBZA3ub4u
5/WTNommKplYcElchreGPBfUF46YUL/I5pe+JB99EclgE3YhTXnjQMg+tfsHoRgA
uVdO0rgKMRIIPYuxX/PxiULqrTc1LLo4SkoR4HBo2qXAEwfPOilqttSd8mrnNRn8
OdG63QLYuU07HQRuoxP19mp+GlFuujKPsz32oP0OaLedhfP6xi9MM8rhYzAKNvib
xKT1sIn4T4lwjWzfu04wFJzE5Mo6iaCrWl1HTpM1jj68mYI+ZGKBurDAapnhoeqQ
39X4ST3vQvCMEfmPKSUrGc0kozf7sXajt7GqcF1DpMuqo4xlUQsnul80RIj9EEaS
SHbh/A3X4ry5nPOKfWn3ErZ1CmKGqTW7EnXCmVyipi4Evp2QcvMzuy6qRi7yAjFT
DYvxKVb/JtRYCtQulCVht1phiTvsvUXfcl02TSzz95jAdWGUfzJHyWaQ5xB0B1sQ
54D3cxx/YpGdUeR8FYOcIjRKRFeaT1mlvOkCUJnOuba66eEv6QbF+bozy3pS9/41
e2oF6kFPIESs/O9HDvQrs6G/+dXeyn9rn7AwvFHaIvVH5UHXW0iNsXi1ao7u1iA+
b45bF2nupz24oT4eRmukQp7lsc54P1tZ0UcqSrObFrGcpRy6M6KONgfmi4TCk9kc
Yz4c+8FyOWbqIV0fxG6c0rTSiFVYssK7a9wkdPmpEyaqfL536yI73reJ6Q5aY3m3
BUzlhODmZhbHlJu+sq3jND9vTAQryXEoXXQdEe4w7Z5e58eiwfxF6qMea1S1KZbN
LyfGm0p2s7KvF81GPcIjOCZcHpDMBpYtzJPLSxhQDKIa8mncT8wQYkDHIw5u58MU
v3Vh+3k3VZQ2U6D23crI94hZWHbWPg+vs4GW0h/C7ZMGEQ99+JRKgOP96Dia+ZbC
ntIsG56BwA8yBdl4sHjG/RhSDDcBkymJSwTuFNxGKyJW+lM3CxqGS8in3mI4afH3
Ojb3yzGkgmDJ+eAlOHOrTKXp+3cUBanaco9D3z5Dhi0KMlUIoa8IG5bicY2xJ7dl
em8PgEVuQdFUzTsBcsgo7Y/1ThZDXxPVFJniLwllgmbdHHAA5I0JI+i1haJFQS1X
POaT3PZagjY6rE9F45IF0wXMe8QiTBqh/jw9Io1uQH2A0Y/GtlFuJG1tAMen0y6I
UgfVW0xgl4DPB+U2maLmTAA/QR+s3m9UbdVASbgM07n9vabgqOd3eu+f1KbK7SdP
4S1MW1YQRBcxcEIgvyQyqFIfeR/YJN9XD/7w0QnUmLzx6TOzYVQ0mmWVspf5KCa+
THvV4PmOuklUPgXQXrjAruMqlmFJXOJKFT44ORoQlTabbKyktHFCDpRqvVI1Lcw/
/Ys6+FkF4O2xAruDPgTCGG2zd43Yv0fzeINqTKCx/qPt0SVrcnVzXW1kHG3Z91/d
cQdPHi5u/o8oNC379p+3ZKL3hOBEIn3Pqwd/yQGAGHR4ECoNCsKV49bjSr1UwJ9t
2ntN+QYXVUFQ4afKSC36lu3qu0HgdhPu8v2DIGZl25YmGo0iBhdYLN2daIb2e+Qn
taCzvB9arJmvlVKGOQC5iCEc75MnTCsYkMwvLIJeN5Zt0CAbfmZWB1zAHhDsV8Hy
lNDZJugHwLuTvLKDFkjNG+J/a8OnCTTej6Xrp7CXXH3AR/g+YUfA9kePbdZZ15SV
ZokQd6zaIhTt/fzWNcCtBrRI9PsX0Pqwcp5ohQ8IehYnJ4rsS0inTyC4RHP3drtw
dw2Y1MhYu0gnhb8tmMwa11v+ffpkVmCv95IkYfVeP+BB74G+nGXpyVz7ynTZ46UU
1iibX8ngtd76u/7hu8H7TrX3/bcRgrFVQpOVplG65esiVfMv80279Rm1HJhPSdtL
qRvPSpG1DOXpyCdAKCp0XmK2RReu3NWXbg+ud0tWc6WfU7NreZ3FgQNXe7lHBLDx
+ZIEvJ4KoWlun0MsSMyxyQ3gHctiBu7zOHNQyK2APkJm7ppGg/7iFmB6Rdcjrk9C
bzSOuDs0AdbDtEVyf3AVsN4gXfW+0lPoUPipMf+B9Toxpo0fDtoYWeVVS0rhDQJd
ilRLGloetu+jZ2U/5s08yuugCn18at+x4HilYbnmHqjPh4S7jCbQ3PhjGx4XMPPv
GQ42JQXMO16lZi6vk+an6Sh0Eu1Lzk6xBh16a6wpS6mrF4N3Rk4qAKR6dNR/33yL
bgIQ9oCIgUMb1d2jWem1LdUZWc5m3DBaRnqdutl0WIT4mAnUg3wOFDBptLlk+Wm3
2xBi4MPtsymFasCx1kELqwsqnEknT8U7ZZWDdhc6Isj8OXa8cmXF7Vns36mJe/r1
PUf+kgTtPm83hXUH3NHKquBPAtVhITXwFe3GTQ78qNdR+Jt/SQQLZDYtpi2mmAhD
SY7XfGqL06ipKtq81mwP1TkCmDZarDtWqdByKVPBoXW/ZJNbooVGF4Z4U4bxq5gj
k3KfxojHHXuDCgXSveigHf95W0bzHmGRS1XR21cJb09R0WxlIsuSzii8fsx88rMT
0rDi0JzIZbWoQSBY7hR+qMfRYG5umGc32qYmk3h4BzgmlphMbyfh+RHqp2/YntdD
j23u7E6ci+SliahzoDngzUVMAY4ll+sdEReEd3uts/fS7siQLXxItKq6QGj6lB6D
DVHc9fOPGihDjJKxxsZuFIBC19Gz2tmsLsm/1xho26BR7OwesiLLlfe4352SEE/G
QlxnJjjjdZbjysClf4FH+wRyGuaJLbvOUq4Jrm5vPM3H4tFSr/UaiCQ64G4Jq5DV
epk5xOdmfqLsQ2rfyBJ4cjzKnIKTG9TbWW6NNd3o8L+5rMB6taKTQkZCvEpux8mF
5VUUwLc/p4Pv9HJmHyHYlu7W6rPXx1Box3hduzvRwDXfM0RnemSIkkVFcJgCBPrY
/QJ7GPQeEDMRbdBtOSIGCoa39RXdwf7PRf8TweNu7nqlzGB29iOUIsVwUqHKklEl
tXW4p6BaAc3AHg853szErdXpDypcM33igvlacvQlo1j0IoB3vGKuL7pUwu+dg0B6
ruLI1/RtC7Ry8tZDNbw8Gairg0mmRuESDfc8SlSlt8vJJihY9EGcy2DuTB9EcCWt
wrc7YztqZq7WqG7zFmXBdRl5HvL7jPkJ6kpIDCGWpLLueEKZn73sBDbi31jenaFm
5CVhVEUMhtbtMzQbkxNQ/FJIuKtuBZK9D9WaVB6sEaRpzt8QSQaVKEYZxpmQqWyR
WKQ8PsV8N+1qxgFeVIkq8sOsWD7ZO//c/+dX/gGVoju1epYSFFNNiDZixPYJRtJK
uWH+U0rF0iJkBaZr4TutvjyoQcl2ElmnTK6co/6wBFuRYNj5AAGe3nl7LwbXTfuH
dBA9bM9qBlBqObLRzVURkvchJ+QOIPbvhFo4xXT28XwUnYrgabkeP89kVwUUwAUs
Az/W9ge/TPVMcyFzF8183US/f50Sn4adErW6lV/ENceWrmh+XtC6gYj9a5fhYTVO
KB6FxqtL6PQMQkOP9ED+ULCELRG06rSTGbxwttjC+lbAstzSwqb7D2lnggfuoIWH
5DfjTVWcSKh4JDp7XjREREeA1avXKR71IjSv6R5RNiGMFKlinq7ppJhg5JyMoK41
e5SsLjUezdbQtrZxUwAEl/nkVbKgIHAJ7EMsAVQqrzoN2wz4nfysav+GBeiHg62A
ddXV7TIJSqPbgTiQzO38OXjIXwYj1MZlhU8R4QIyjPQwkzc200QN80FB18tfJS9E
jdsLY7SJjmaFrpPuM7JOvoMVLJw0bAmmc1EAGF0jNDITxQ8MnLPEDkp1fHRFYSMH
LV+imKj7lOQGYoP1GNYmqKIJCHqMy2CbGw01noyu2XYdd3+1ssvX0QVuUvgKG9X5
sAhC3PgZZSa45pQySi09KYm8ciE7ms7OF12ZALXZHpDvN2Yv5yrS9Y8+7Td1/VY6
gYhSWP0aDFDbbw0bxU+UgEvfeDGsfgzEkC9lEkIH7fZ8d07hR2T6JrXO/NPY+Aym
rqqOp0aTo1HVyvPiIcnRDNJC9UFaUsW7ETgnpur5CmWcZyu4odqeOwW3i/sW/dhs
boUS81o2jDwx+c83KgrdLvFX/KkTw0kRQYKjz6Wa94ZVUaWE+aTv9slGhqnQaD4v
2HiceTHYw19sqDWTYzTkF7wA9yG/8SnHziKKiXac4mGuwRdCzaGxNM3isHoiqmCK
egWGBNmuTwNndHlTFsO5JI/vP1ognRc/62odRV47FKk+nkmVdDxLsI1R5ZMo3ft8
31AxFG2aVtrWry01vZLv8bU6kHpqE1gpZu/JZH6t2QHmy/pNq4YXJSXPCLbvy4vk
6McRSjIGgax/j78Kmg1kDFEyD9x33p1WQxQy5a314oy41dzolMWX0s9nm6MdavUA
iCDscOLcsrZfSJzZKwliz9OvJNIUlntkKYmEeCump2EbLGTdcDXM4VmPftGE0sy+
U0DfrlN6ocfQalksB31HbWzRlcqHHfD27y4RZUp8pde//3XIK1+XsZzAra24hyHX
wXcV236GlqLxwR4blBtSCU8CW6NlQjGwZCvdHahxZzJOITHsubjbupcRIXZINQTq
gtCH+1/B0bkq1WLpZ/e7CuX73fvMAJgMvDWeG8XlD9J7RIhK9Dzcgzl7aEnIkWBY
r+aR4YCjWo5wL1zlU/OZhec6uzUmm3ERXSpvxjQePCaohue2zIvKFlTnFWFS0PbO
uEL+isLUOmnaa+Wvr2U3ztR1RyqdvCWhRNap/JtQfbFWDeJcMdwVlV1KOv1/TV0N
jpLzmWdX3iALOVLJQoJfgKyW0/2xrcYwDlECond/6tc4lGJbNL5Rl+51WI6dLBUI
oFbzRuDeVL8uDcpOeg2uCM561tS8uu0+xK8MdzCnPE+jz1BaIkjbyf86I9DwDWX6
kWgHlMueNF2m67/XZFuC0m+2xeKPFwcDlblM2P+6o+YantyE+n+GmagiIWgaoM63
s6sPdD/NDQXOjsbdYgRBuCcKY9XDXu0IkQeWB0V4j+6OtaIfNjkYT01/wN6RYEwI
YQsADwgOhePv1gxxg+ap1flhkLWgRY44tFF0VOH3nnsAOdQKDZ0Mkjr/XaTnW52q
Svg+diWUXT6tE++da16AbB0FQ3M19KPvPm65QKwjp6CZAVqW8huKQ9XJe6x6IeFD
jbq39s79k4CqYx4FtmiTwugf20bo+rKT0KTwzVuhS4Jo+Ez8duAZ0CQhgiFzWCBD
mVUWU9h/Yti8QKoRSJfWMQjwjAohW4pAM66blyN3EmHtskz/qwjryJ6lJ5qwJC3L
5Q68FH5U0PBWouW9GzPRqKk3FJ22poapwL+5HCHQ/udWcRVs/XMOl+Cz5dmvbclf
mxApkhaAcaHqxL2eZ1YEkGFVlJAPye1hlcHc+6DwPS4SuqjWc+SQuQuqKxQsUvwd
qxd12aLW51zhc2pbPi816bhEKLf5MRyynz6Kka5auC0XXi/ecBNJwzXAngwDp7FF
xAsM3rs3YAS9gM821ssmAgWpvtoGa2LxoCv3p9wSFLFugpWVKNM4iBsgUeYYik9a
5d6P+RcaBPlOs986n+LmACvRdZ+1HgVqrgQSal9AGLjFqeqk5xqiNrhfSZShIeFo
Gdn78J62bSgltTXNmK9kkYzgI/u9dseY6sTncw16KCOUj7uWL2Fw2Ph7844JY0kN
uucPwXYQYlIgU0OjSNNV7LBGVCwALF9h8AbM95YjSL96oMZLV25NYiqlXU05UCKx
p0ykcjSm0B2DeHOciBaiiYlCQxuGsul+gxMAU7CC1rc115hPjWAcm6SD3F9UmSbb
Led7S17X8AlTlDpgu4FJivlUrBXYDBs4bE3KKoc6rIsM0U2mBw6UVXFlhiY59aIr
LKqGAifCZDP655ivN7HMd9lhZP4XlG0bhMAS6BLDbNsuGRm3MMERDmJkw2ILTjd0
AYPJF9pggt3udmkPrZLuEqXk8nWomClmzi2T3WBYN0BX1tpP6sCvFdeskKJOqPBy
UfxNLt6mb28DIuwCijoaDqhAOg9UTjEvSEEdh2RQDY7uBSL954ln1p8cm64tsuNY
IihAONEHCRXLBGQoMv5CB3RYDU9tp63oXLBXBgE7aSMOWNEVKpUERAVqfhdnuNpv
6KD1noV83PxYqjKhf4eD4GUmLwZx6uXq3ElISU1gkDDd+XrECGIclkPLq0cs98ok
640bWykTist3fSQhkmCdwrneEtk+Vvz3MFhOYjgEiex3BOI5w9Dx7LJAyefHm8bj
ro79M8B5b7Hc4jp0DrW+/bENY9wnC2F6hewmRjGIW/VHsr/z9SEcYRQDst/ZbgKb
esFXC4oB6jjwUeYC4uPewva2sVrezX9RQHuMynpKRyqU/J/GRlKaFe5eXmyt/uwi
YfA7hBzFyM8qS/qiMJ91w7BCLOrAJEfBiP+p1GvCVAT76W4xf61oTfMBtGJ55Ixe
EtjTGnwZ4R5Tn1Ts2Z1sIuA6cD/B42VtJH15iWVYCF68xovZ9+VatgPyvXIMrZOr
G/HFBK2OZYXcNUrU3wAQYSA2jD0G8rOpxiLW4DNRmgMKGZz/nlc0m1UmXEbRcuaB
+EtEPhv21M0QCOaVREIvESYDDm0ZS6CiWjtBuCyApgNMiEc3Z4v95MRGYkbuyalG
F48+1JZkrz0kdrgjcl377U8o5sULD/sWP3aA9J9vvD8rygCK01nsbidppcLVpKtq
zgU4r5PA6W2sMWnvsxn1MQakuuEkK6tYBowvY46Hxc2hydOg8I5udpADYcYeP18e
+p82b2JpkoeQW/jQs9k8RQGcHlvtgPpwys6shUgoYL9mOIuF2/oX/vrhrQhG4hhI
B6WddrK8kueM7IcdOoVD84awZKBpdYoKMldzAbwUlNpVWxDKB94ZrZu7TlOM9wnE
2NCB5nH+4iKHaz98peAwmK/kQ4YmiqBEdrTfxNuESSQg2Y0i/uva0NDk1ohsF2uU
DslFA/kB4W91iVIPVt4eictOc9guf9Z5iHkgQze2lZRirF19iT+KS306QhC9V4hP
5EscxrT9RsSK1xxDDnJqT5HEHih8REE12Lh/30sdFJn2byt/lC9RLe3VYf6EZlUM
y6B5EtohQ3UCkWebLE1ypW3T/gh+tkIkG2UBszBBs8R9h9r9/pn/WLG6OT0HgxLX
rqxaYNenvsFPK/LGxpyGZELesvOFeitbms8ngOrLzXsPjvSBAWryMpInqUksvYpo
lOkmn2mUzp1Dx5cOVqjV+QWK9o4KnirdrtzmFg3YyXnG27OkkCKc0xigTfMkxMO2
r3NZCUJLbqi3U0NKiocBL+/LDMNLdOaLpFiYMI5qt+KPDKjgyBtk0zzBymElKDHB
S+UsDFJVA/meJ8wT67apfWCChnkwHIc/sgq8PhIpR1PQzY6cyPhoct8JmRqIGY2K
OQBckNL2UgBOXQwF+0jNdoC5NEA8vTtGkytI1Pw+QHKpPfxI8IfRP5k7m42S1uIj
q2uCc7na819wRUHI4Ilc+j3PEdTr3WylgqflQqNo9VU23eaZVW1ysAXEMt8EhgsY
U1WcF3JARuWPvMmNcZ/sWfCzO4BcIKuj+tTSeWBoSVD04xT4eMMMsOIUzI5czZYv
SzCtnKJBSU4l+SYOg1EevUG7dkuyQi8/Q/H/wtc3/Uv0Dtm+5J9p0+aHWZ3M4wLz
nKjJ94L8fkqSJb4V9YK/ByAELlkkKGshu1yaq57KihLsBwmIQTOTvppP9KTE3EbU
eaV6km2F3zgx7V0eE15dYUemcteBzl2f/aHiVC4zi8kBhcQ1Qrzf/v/dYizpblSo
5k8BVYTAtq8Z/9GfneGu5gcdZxdAP6mDJ38mXzgx27bydhi45X/oJ94rs1vBpxTB
Lf/9p8zauavT3Ji4ehrIS0cI990d5e2u1bAbyBWzZ5oNtadNDCL98bJ6xE0MjlcH
ySMj7yMDIRVIVrvQ9M5aTiIlrt02ltsvpxRsqKq2zVG3lOHQmHDamBzas0COdDe/
iPqDv5RnztuSgyjrGOZxYVux3aZlaKpxwrmBY8bjXIfsewM2zhxfAAE0D524SJmb
W4HB1CjYlNf9fGICy7sEOEIoS+5nwy+a5xzP0kD8ZLArmOrTk4U9U0dsN6v1Lak7
MUfB2eH8BaaYs844owm29YEuhR5Fe9A+kYmL9XLWTWopxUQ2soWHlMBwjKVQseph
0HLWyCDM9iA+gGJQ2VqMbCaZVngONUd2r+FuF1hy5btK+bYbth2qK3MK+Sc0J/os
wXmYv8LzKziTEOPsL0ZZbuMG506/P6C4SMOdIDhQH4iM63OVBnH4OnUcUJFJVDnp
cb+G9/At1sDodPFkvLHkYpu5lJX83HDxHBJOiE9fm90gLeRuLIL9h4OWPsMK+q9c
a7Oi/KV9QdWoUEBtJIpDEgogqnuvFU/BAtep8DYlNHsml3WquCSa9673NUUcOu4Q
UpTcaM3S/nzwErK3RecLIvUyQlwfk4CPYYskzA12JcA0pOrLX3bwDESV77VaO0MW
oAa61YiUaj/AngG1QDe/cdCzMd5NtiaZ5zE7qXYqu/ywIy+REYk+6OEYW3MV2TGu
polhyxXKfDexVKJ/dXuJRAQUlCjnFvj6tfAmdo9L9l0ms3aWxs/Y0vaXMDgAwLhL
X3C7KQ+QCqDPhV2dbNvG508+irP/cLrNGg7b9yQ9bSNu2pX4pgjcENEcO4BcbzYJ
5VB50CUxi3aNBjyYnfe8qcdbYX94vpT74z4OehUEE5RCRvuULSihWHw0TkZz2PmW
D0KMckPWT2jfQcmC+nClqxn2NBNQ+vtFaG4gKj3kLGYJF/2H6NjNCZZdQv8G5jer
uq5LyXbS4oAXna+dJHHTXbcLgAxQcsx0IOH5tF1lYvlO5XKODx+Wy340nH5USdmT
fqxoHKbp1mYzgLG5OorogHgRp04FeYZPahICSeGdlpIvK0WLPkgXV0TpAqBR2EAJ
jM/BjZQtl1PjGwEsB67pWMr412XUSGiqPE7syhQRqHKWBy9vM3G+u97Hpj+NTLr6
VKKIyXec933NXo6Mrrx1/K/y4Ul/DJI8g81/75EI30wzTBcs8xsLnM7bsupnkH/o
o+H41LoL8u4xhS02t19LKvRhpIyDlBdPg5fiAXH9ceoDIZv9/SjbsJplLDbRMopv
KZ3Ereh6N26UULKLonBnbEJHHBWXDsk6qZ0ULQ+Ey0xPHeAy4f9825wT1rJnonZq
AZzH2wjKybNh4e2ZnwaHcIcmX1sVMkmbRSW+vgKOa40nSoOe8/LDDUj2c6aiChqp
tEMpSLzsiPpeEPuYZ7EHwJLn2RA9RrOltakQGERo3jeXyhXcEVxQqjePhMwRLCMm
MEx7s3pTLPBiGFHlmyVh8eyYULAcJzZDCasx12GvsMVaYwIz5xWNcHHNLkIxCcpD
eNkT7tcytV1pxjYitN3bKebDsUBaz/RTvPiUtBbzWpQXQt5tmjRj4vERQJRkxxUU
U7vEYftXLj+txMZDsCJ4x3al5wFp5SpSI9yxK+M2mDPUaIY3DwnbY0hdczRHSLn3
cnlKLK1EB/JuF2uCGXguPEGA4QeC9hYRqNrcYwMISbEPvOXLEc+slLOHjF5vh7Ub
fCWmkgQg0r9DQ4RG2goXYLE78QsblL0gry9gHz25tRzCsSQ2U7S/FLYk4SiZ7I+f
TeiuneUSFGja8CANftVOiKkUW8B0o+fQ54lrATgcpm+WjwQ78A5on5AY7+xiKzG3
t1TzFFWBpOWJqv/pkeHbbXMDkcUskEGMKksc2FfgEOC/7KAyVCIJr7xx3iN3c+xr
/IMmNiRclHheIRmc9041GuT68JV3k3VIkpHwHtCEcoUzCjwwn4BL9LzvYCYmsos5
v8lAJLKJjfrIlh4wWrUztnYCFBG5N64jgMSLidwBFcmg71Dg1QcPiYm1TVaCi7w9
iRbMqQLusvP31YvFopJDL8HiSwKhMxy8l8QaRia9bh6UnOlLbdjDJE2/ojAcO+jA
Oc/Gabo0uNw2dg5YdSOOH8zI/Vb5E0VhMxjaLOdZzIro9jPtEVuA8rrho4SrO9rq
xZyZDDV76waGbjPAKjgt14zVNURFwpy9dRBvnUhxlsoLqIeUMjOKrZkvg5HeeZtm
kQECy+2FeA0jJm/bD2u6HfONLipkvRuS2orQU4I+fXSRuwMWiTnHgmxOHIArMqNx
bHJCWplo7BU4fBg46axy+jya0ts24yyNpvALENfJUOf6+ELxRDZQgsPK6qn1a6wJ
YaImsgg0c3QpJffFt1kyO3Pgpmde4Ub4SgZiMqLEYDp4vLC6Z8/UtQ4Uooetp/Ql
+Blr13K212ePwEMC+Cd3m0lUibA+AcOo45ABV0XR6QWHSVXFtpQdcaUeoK07YSzc
nu9iBKnZYQfZrvZt5/S7hL4TKnEEaY9CiJ2OWRPcPyocS0qPO4uqw6PJJEBAe1VP
I2se4o2/xreoQ5AvWpqdHTAgNAguCiVT5YUu5vmnQesvVDaASSCoDoODyirVAuyY
sQdi4BJuW12diOWBFZmpWAxe5ig4R0Ws9y29S9nou1wspdlQvZ4bDZi1EpXOdsx0
cgAC5WyRe0pcUGYf5zp3HjU5rXpvTSrHvRCabcVh2t2A9rNE+gC0z+Q7jfaJ7lCq
Xiyx+IKnCYwN2+qsEFR9vVE7oBnF28h2kOT57l/kTKQPt8rLWkAkEgt9or/v6GKJ
Ft/YH3+cHBraBbgbQEi1HcwiAoY47njuVi4gb8WXV8l4t+/frXK/U70rPBFm5jaS
VDQ20Z55MlGOc2UO0YVTWG/hvhpb2IYSshjbW+V+QuLTJzMdZdydAMmcXWgVmO4s
+UMDpVVuZFzDy563VwfVAcx+FQbQGJQgy4VgVzjD2+sbpJt0cuYfmlY3Ed8AmAb1
ZDRxydw9PqaGftLOud5KSRh08XlXfmEns8LBIWFKoYcfwEnLg0cAdGJLLHD44w9j
4p2IRG7oPe7MkBV/ff8IyxO+k5/CVTzI780FKjpWfO2LMLC0WaBn4Vc9OOGWfdCz
7tuiwB4yzQlICzHAxtaAXPv8TkZhtHQlfGLQkeEroASUkKlKmSAWlKqSgFTTm8pw
5elW2mWw5AOl8UIkG22xHVLooXZeJgiioMZGGPK3QasEvlXrekhOsmd1PJeI5tAl
SveSn/2OTCKuECo6ac4ercVLWe4gpuJ8+8yx3F4U8DnLfD8fTE9mMTL3WYq9z5fL
FA0ZJ1WT3Ayblndw0SMRrTPJ31ONFZ046SsbrsYIwNsK8ZECEniMrKtpmwM+DYLg
yLnbDQmSVHvr+ZZcRdH52GYD5L/NOZci0C7jyuMxbxmIoRXws5EDbLTU4CKDQtU0
2iixYZDOpYqr4vb/ajUKOhb48mB2RStAnlEirIcRNTEqOp7NX5f+IgWcneNVxYcS
wrapuxnlMzQ84EO7H5qG8WOG6Z9HeoF7oIWT0qWId0mbGBBXegIkJVY3rbbMbWcc
s6MEgXC1kInjKFKLpOFXt6gAxlz859LEwDpCE9n3VU1baeaG9yuVNxQJatPJPOkx
MED/MSoKOW3VHfjCQR/Zcs7qAoAIG11ApyNJnjH4vsYQgkUFTMom5hY2oPjfZF2a
0hIODMhPxxuecaHmiHD8TRENzJMvGmQY613fRMf6C7hEbUPPe3DrsEZgFcG2VjMb
FSfCaBIKoZqFSrLMAnK/7fOqHCo/C+U89lT1dYUOiROYgCt+XMyLuf9xgC5t4A0a
jULeWMPNXQW3RhekobSzRfp0m0HtvNciJqsUQ0r0xoEg3bl+7shtjZI3bFaFDvIX
xtkwbjR48GXWsviGHVvJjMVOntS9zeJctqJJ9ahcC/N0G8sEDFV9EpbL3Zt5/vhb
sksTLg3/BkekkhVpz4aVjauF9HDlLPxxHkRNw2hB6ztEzCsFkHIBFeqVWA0uEHxV
o8EFC+os2jPosJ5hBT/nquCZ4PVMzqvMbAwUoIZCLSb95Hgmeh2mcX/08Hayt7OS
Yf5rMG09CPS8CE0ugWjJyQ4LZutZlbl6qHym9s8Ny5p/Li1kxWl3nt+zg/YA655q
Wi51aNV92OmDWjRsMn26PkYE4/C5glx7SAomxDTF1oEx5lAIuLMH06iEEAgpM240
0U57hwkV9LNPBkHOzHnZ3LFrDsYv4IdjCaFAKdZXWhSkjwUbg2ap5Rmtxx8QSUD3
pWi7NcT7QTWD58yoAdQtHqToZUl4akSVYZjRB1dY84eTe7hnfLmxflePT4XGz6Bk
j3HGJY9xgo4c5zsys5+1/4Wovao9AYW7hmkYSMRy488+yUqmlRFIJzP5mtqLSEbu
rKqk3OypaoF9+ub8RubJOOp/b1lO4v4QfJn2zXMEGYcLfuPK1xPsg0u1U4zDAOw+
pNKQ/OUj5+6SQULqh+eVMjOsZWVEdImBZp9/9rdsL8TclQuGdSrZF+ioKqBaX7Bb
moS4di+sUZb8xHAGCJVVDYIXDtP+cTcVvSWq74RmNPvvL7MQ6f/hgdupybmmDRtm
MFmWaNce4YDcaStv/KgrsC0x3JB2Fq/Ct57aSupsMhidnJDnLoru3lZw40sIDBhq
M05RFg4kqZIrVZTK9dJLokE0dnfq0IMX1MVfCfGthDh45Y68tKS6dFxMFWwvYTE/
daq/0q5YSD64BvaK+1DNq7SCfSB4uXhV8AlQU3jgkTvUqH2cpO1X4MHEfs2RfKwV
fI4jZ7kBjcW3qabMW3AYE98jBh+OAlILo970xlXYc+16e4klPYCa3Qu41/Caa9JK
wSiDok1v+xUBgOaUvMkt0q0EEnnOH99vUvzOShHnKMPmnDfQO0PPqKyazBAJgMlm
4t2KIQ2C1scY7oW6iUxDYbwF0NJngQ0qHJpJMm+vtBqJ0ULPcXkXAUSNTWdTXLL4
HNz9U+UYdTYm/KaTj8Y6SMGgBNzkW9qz7gN11nKSm7t9MdwGG8RN5+RwGfLIRIJ8
5+JT+EJTAdaNWM2rVqSt2hK9m7wYoAfZoil/MCTSF2NuB/m9HEDS1Lrnz454Dsr6
VpFhbh9Dr9soegKlSYwQ8lc8zF1Tb52IpHEob5tT6yLOXn7AQ/BJWC/e+JSj5+i8
Fss3NwsdTG7easOIu5TN9nNvEoAvUGoZYY7in6jbbqT8tp81BtGSN/ccAqe4LIkE
J67nQAY4QfcO0/If1fMdkfQTlo0WVOsNS+ZFvZrZE+dKt5vplBw3bDsgvSYaFqsf
H5k/L+ovHrOj+tWsktwKnlPcQk0AXsDetfazYsdm/+oC7HcnmLo90J1RWua5aARE
5At+XkIgHwyqKCR/ufLxSbj3Dq8BF3YxJuoorBLtA1Cg+5yGhe0KnCcNKdYP7IvC
QYa0hv0ZmPTK9TFpoxrCaVPeSNEFutME5pYv7hHTC0Vfh8N9LVRLCbkkPQIc5Wq5
OA1C4Dax1uMH5H50R+QC5RTAATV0s3ujBxy8dlf6kW6v2Puksyc9PRvhOBvg+M1+
lhYfj3nN9z8W2/3Z3C97iymqV1kA57dfw1IVxNhBzX/QxNFrZLnJNDqJpwHnk6S3
DiM5UGqkWu4ASLdFD4OSzf5DjyF+TpEx+tXQ5DOlFmGWxDQYUGIujU6zdSy7Fthd
sbLpfvvgVcotDl/MMNEz4SiPrcLApngSzRZ1eQnhB8ePkrBsH3hY7XRSlGcHE5C1
QK09jQj0PcCWXBNEQ08OsFdp6QqlU7dFclSdBiW2HH2qb6vNT2lEMAQX6cLKqeEE
UuX6+9Y4eLO0vv62CRuv/u1L5E9BHGQi1NwYuwpKpnja0gwCSnObO0usKrp4uiTD
IXMi/fXtZaWLROQ1L2QiPBv5gV/5K3MB1rIFAJRgB6V0bFnxj2CA22Hx9G4qVNh8
ASF9WVta0Ih+EL2AQH1RorPNP88ASxapvS6CiHD+/6VQxacpQtuJpJVVBO23Jene
TySo/4lk671JQSPlqHe538YjNolSfCgOB8EIWMVzUN1W/GaFmAylms3hA17rHD9S
AKvi0WTbV/ljwgpMf8S+F/458KdG1mkHu8QIPiGNoJiIRL4pYkwPBvMYHuamagfq
kFzQcNsJXaNw//n0LOzmjO5+WOXiGaFda+fSn1KnE65z6//cYylut6DWTVx1SP6K
Y1Inkirj9SxqzX/zG1VOeGb9ACsHNpq79Pzr7hdmEzpVj1T9VmDRiB82jle7l1gi
XKU7f37a4Elc3qWHquYgh4x15Auobzl4cF+Jwo26GlHbwlqhQ2W5kj8DnEdUzbn0
5APOX2zW6h73g/9KwoLQShm2mEyqzOOI61aLo7e/h9L65LzKbh6/wNrtEhWLtorg
phJkiicgXjNf/OUc0QH0g9bYfPzxXkVj5HdQ+pjMSqohS15Np6C/4Xjmn8eBx5G8
o2oUON3YlFcjOpTGSA+Cvuy8wsSTg5uF2txD42Iz2b015lkhIP5qEk+CqNfK/fqb
9n/iediamBNERUrpXG1ZjxBXmPjgfCGL7x6d4dyYll9pzP+ieBtD2YVv9FTodw8y
MYn8mo/WxWSvLR4ITyiR8RiHoYWg9dm9n5a1IMawLBatqyhVKkQ6YQbz5DMocY6X
z25TAmGsa3EncDW2EN6rLUCioLeBx2iq74KQFHoU+Nm84T7vVTAStt9sKzCSDJcp
vhRFUMes9hbUXtqS+tl2fST5ZDEL2YuD5bPwUlyp+Z7qkLglE7W71UFx4FK1SaGa
2m3bZP9MKwgH168t4tShSy1SRZOD7WgXHePchwbStVmMND4ySDmcgHXWBl8e6zWj
dMAm/S+pa09FDP3ymUdFrIJt5kyYzKeMln4JCc5urwiVPztgDiRQNqZ0mU+2okns
/ISWJ/dDZiWNJGxkEeAdm3DnIvqQ4biSi5jTLg7AupPnaNHFJuxsdT+X+Zd6s/qx
RURanZXKT739lBFtwQTAV6FrTl5aWIh/CYZO3mWliFSmNPzYmDysM676gA+V0SHH
AZbbcvHrkWdhyjD3iZP4RHKddZMbu693dunsJQ68tYHGtqg+fCDPxr9VYG/xlJKX
AjbLJbvqy1kS8O9fLQuA2FygMsiURqY1GTXx5Vnrq05MgpVhRBnzuywvVj2XFPEa
iM3/VQWF8XVXPP7sJzakhBqX2vUvGzdqCDw2tmJPbcd8rhkjw58zlP5gUn4bssUs
OBUvU1LnAxE9E3lQ4uMC34v7FJmqqkCV3hVeuOqMA9emLNRID0VTR9rp54OF8gvg
/reOr8RXfBpjcS5IeuEo6zlcodySjoEtmzEArqqbxLKTmQYEBpSbEuY0zeogiFe6
Y0UYxZSgtmWy/uVRSGh9kxn0purCitHf/fWoAYuHsEZAcCV+dlYHwFg5gX0fFmtY
8JUr42Ta8VyE0EsgzJxwBQSN1TV+AiiCV0yOhRVDPxI5kihsY493sfrowz/WXgNH
57ToDtmqeQSSbGBsbdbP0Nx270rolkjhtz3kxM+weVPw/PqSgN1ALXPFoc2W21e7
xnfKu/YXXhoMHQxOVszN0I8iQIGLVWMTzkOcry6bMB6JmXPO1SEtRvYDr018KoY4
e0XiaXwdcqimJLkoOwHecWbYUXFco4pU0XngHN5LFuIa7OzxWpwphfIuxRgvTPuV
ypvKWgc/yNaXehDLPZCcKY4HvqtctQxd17xtvKp2jK77Ig3URD1wWBPwgR+ea32i
WVS21A/pW+dXFR8gDrkQeaCuhF9YFyQTeNoXr6IiutuiH8lkd0p6A1+WfR+lAoXn
nAlsijO+aOcKdakLSw+Dr+OTSujEl6KqZXcNp6Dzo1tOmHzC7uAr+zwCZPw0eMPu
HhNSYjXWg6V4yCp5tUfXERXvqpd3T9VZf3ZV/z7XWKWondCTe3WOQz5dO7hj3OMk
HpnMCVUCN6zSeqEkqzXNw3ZKx6zFoMqeeA67ojoYwXKY2x3eJJvXImar2O8XSWDl
ZEpRwkuYVyoBRVUnRnCBwyBwnNBDy1P7Ryt6En12Tx60YTGlvROHoLYY5xfMDUIl
K7i+rn80Re1n/3qAYzBUbKYrF8+ncpraeqTvlni8u/E4Kcbh0clmYTKqAEeMElqF
vS0nedbZlZqr+g1KI+k5bLBobfdV4X9I/LtzTxz6H7xzlxB6Qml0aaXq7aomi1WE
fmlMwBKWCNJ9n124/neZAIhltvdVpzHeYxETuB1uhdP4noVY+hOSMDR+bV4aO0Ap
67Bnt6OIq8Pp4QH/gLYxymg8Yipz9DYF5ZZdT3V2uh6dAYfBncUC+Bo/xk3PtN9p
9gZTEROKrCSnVbaIxQmdTIH0fesg7yY2j3jKoT/1+NGUEKSQnzmDeURf6zRGGb5Y
huQBgQ01SM2U36BRXI6iRpmGCKqdIb4k8EnL6umCpSuhJUV5Zw/MfSMhntBpwfsM
W4sdocUpLflbopxM3h5RGykqDmttxOCELsYFzLmOCsBYbGWJb9z3mJpLTtdrqNsG
8QgSfKEJaX+i28oV+3pTYCMwLgDyFcNX//ivTzhQWhFRPsewnslZ/6Q186XtsDlQ
pwICL1jmiSmNoPq8TaMPbP5ZqBFEnXU8ZnNe+Y1syBJ+t/0GJYc2085/DFYRyaB7
PFqsPL4Y4NGWhfLIAtcb1z0DSJhJNskh5RifzirW4b4saxYW2Fjjhf/cG52BZlUv
pdOrOfbUnKR/nJAFrFc9497rHX+xhJ25j4Nb5o5Qj8j+/jvzbPhwo73ghb6QjuC8
JKEGuApAqnrnjY2cc3NCMci0IoUWvYizbYtdHG4U+U5nBjMFCCvVwjkuwMgj/ufp
IW6IZ/8H3LNgktCvLDqOL929kATrWrpPy0BZfG4M7UpwmA4ejUJ2NhAgMZqyFgPK
0HwzaeZwQrc2GAkh8aV0CeBq6w35qD2kjnVgNYbwVXzY/JkjMUSWYDEIcZEqCuv/
Ldd6e88jzBw6TdQxst3CAUgfRDq/lHXhs+IXLGpkKQO+8wgtdn00PJwqpw5AdXfo
PAt7lG9ldj/WLIcIyEeumNKonRFs/5CvkD+nptcJQRYnoteNnDM/ZZSANVYIYyvS
YejKRo8UjYpuGjJGzQFv6idMn/XTrYGeOwVCPa/L7Hk7snzioK7qyR//SLtG3n1f
N9ZaYRZOj7MScv1GGbFzqM4tnaXhoz1SsH3nhKU8iNerAjf0sXIDbYWDVx2W+sG5
kA1x7c8dyuZi8oL9DOoCiDaM1n6MM7M0iiitbuInlzxMJ8TcwGBh8rsGI71WlBtY
H+EjZceqvxIFA0xkS9SVKvHAAA3sNLpBD0L3U+kUFOXTXgyYKlniquBYCULfp0gJ
/WfyRWfX8j93RqeF+7enIzatfLMmDKDimXPe5qOpiqHMy6YKlPtyyxmg3GOJ4u7i
htQ5uRmplts1nltQN4rJer0EBOWDk6V/6zIHjWEFOy/x/6MpJ6yIRgsYsQMh+cX2
9G1qEXnTbzxQdr/KOncvzwAAG5XGNsT1yvPDITIIusQE+V5lFqa0p49nop0/j8xg
f+2h9IudBPv1ZTc5CbCeleQMuKHulxpQXmtyMP/FswnIOStstkX5NSF/r6nftzQh
MTH4XlA5t6kQxUXKlIDxB13lvJ4uYe0jt5WWZgb5XRrBfSgspp9CuH76ZHfuc7T5
KV2YBTXOwp3ZKPQqGAs2IHXorfKNkj+2rZKgK0pmFZWuDxEGbChBqS6gM7MS/NvE
hObcm7PCKtDte5P4DYCGWTJ8qpitdbf7DOG1tNE9YWB9oJ6Lw+GL7++EYEmnWqHQ
cJOig+A5yrrqMmc6E3dI5rhACHuGquwA6Ar5lo1LcmfQg0jS51LQGt1+O4w60Y8c
rt4uCm7HXoDCP1AbaXwVJO3vh3wCAmiDfwdARusHHv98wbVWfJX9KwxSPIODlecq
8MF+AZ9FEgWwJpipIlEfoqoIx+qKjopvpQqnxxN+JIW3Cmzs1o1iE6kzc74CETd5
YkOMpIBckaEcuPWAP1B8AHt012XkDDEqjckI1wEDX3bXsamDxUQekqfgMy4FSu+V
TEcvx8HKfE16VhxraKJiDti8AzwBtWLSo/xfJhasVFpfnbvL67Jpa+cO6F8dGe8v
M0rlCfZj9H7WsB1ZHXtx7t+95ZSwIWEzX+FQ8hVizi39PDdrG33Hk4YLHxc4Sy6k
x52aLyu71CpHodUbvItEwwWHMWPmROtXkKu/u9me8Jd9JS6HKlQxWUwFRxJE+K7Z
vzOzIRx3fB0wBebjBVki9RjtUtEJLK3ynSzyBVikIYpQxLFnClVFYypsMll+bwd0
5Mf3ytl8LVKpD1xqdxj6lDCqRQIUUCnMEtFBr7qN3gGMbv1gm7xw9goz6jFvEEi6
M9xAnIOT/v/I2jA3tsTn9ewdD2lKeB/LKupfAvgrKLUdTgV33BAcIRATMKWso+KS
nbuGctkoEsJvrrXcXIIwpGYbjrbOcyOeBNdSJEU1Nu5C82woxaenQj9y6vxLHEyl
h3+ek3w3chEVpGA8HoFRE0gvmyGDVvve/AImgJK2M/5MRtCo5h/mM7ka5U8b/3En
dnJjahfIM+Beaj6aeE6DPxzzGItLC1JrCGYddjFtx0iSd+ic/sgWiSMazaEy2L83
rrXtlsNqYtO6epa8cU+Un78DizZ7YfR6p8HFUrLJqmnLAg7JFiM7BW1noozvI7z+
mjCCGVthrtQ5fnHScLeWRVZ4ZvxmwTWLVZgZRZpR2/ERilSFOqtBSwFlmFyFhfHA
gkOuEsrUf9rqPFe1q1Gndty4CAfwxS4lSD1FAgRE3PT4ylCdZ1qjR7g33jzn3qn4
hIGFjzGN/ddhtrQJ+2Ms6vV6AOWcczqe9t1D6Cor1jIMGa35RmzIGfvRkF/dfKiq
MnlP1I9eymKJAMfjBC896Z3iDWoBb8F0Af9NODB4cy8EAAFGmGRvIQvJi9KnkBWQ
/hSLhL8vT9dSmkQImJOKy2GEMEYmklMg3bZ3tA2GFIQ4rJQp9GcEIZcT1WgI2eUr
KrwFk7Y/KMqhqgPCz2MSJqu0OAuhjwNr+xNRC2sKfHvbwFi9J24M0iVE2xCkMntv
U2bsUBEgoViW13seFfxfz9t0KIEvh5nh2v6SZoccBBHCoMK5Rmn9fv5Ho52nXsVJ
Y5eOSS+LvN/susmVzXkqWV0NwLz5c4tbAnKazIZbsNTae2UODyAmkG5haw5yJNyR
KlUWUCDyjOuw5pN0Gt7VmGrEGCkR5qqVGyzlfhIBOThlvPyLZ/AJwt9vIrQUswt5
pnet83VToAVKeguhB7p/aEEFeBhSQczCmUdbdArThu805L/pkQ80RktMYqITdIhH
sNYUk9mRDqxCKUMxbVzh/A9I5JcDuOPJtSRXjTFCYLdPMdvCgZ8Udtv1c+MI/TH5
ZDT35kAa19Vnhz9pF6u0Y5KOCmZYwvkmVkeeA2trxplphrqGl+p+5QkWvS3+wV03
KiDyMzjdLbqW5xfjzH8YPLeiGAAE7piFDZyl9hzA8WurgRDTOZXS1oLYsN9vavMq
oPGw3/P9mXA9XLBpLM/V3t4kkzJ6W+9uDWKJWoIIRj9kxQNKpC4riXfzM6rZDj9q
iWzZtDzlNw9Jnp3Zh5d67Tbu0qA06x/KtqNx/jTZZMhJOCYSKVBRVDYNxT32r9Lv
rXu6hhJaXOlffmcQaAUfA/QPA+BRAvZLQHdtDLbM7tWFdd4LFqqHkNCRBHpTcYGh
007UQJg+EHh/A0/nIYW4NB2pKx8t03Ekat1Fw8w72REzMN88hf5OlIxiew6+h7fu
m12l7h5ordz08EvftZpofxTFbSG2eL40JsnZ5e8ic1nvo5KP2ZDQQiaj5z9NqRkv
JWzJzEtuqIXPR5etUtrL9rb014+F7q1E8g8MrS5OYAj7DrHTI+mxM5kdQchlJtfw
R1LixuFEchzjwuHl/GvfNGtDrR/6/8esfYiCVu77joQIvXx5jvqfofrFeGO1snvg
Ex5MZ9K5QvQ+rZYLNpfTCyC8BrcPwCSnxf9vqk+emMllA2gyiw1KO8BonGgJfEWL
uTsB5v6k5l3MwaP4J4jRooz4s29d4d0Jn9HS+tqlc+naI9g1UMOpxJ3qG9FMRZnw
q4woSRAOhXj4KIOs9kGRcLDRbM9hB8/0H1Ix3zduu8ihe+iGd0jWFwng7cNlfD8X
HHtEcBLaml5yMfpn5x7sHdG8OoVO9bAUC8FA69gWpuNkdGhqYWWaC+vSm6Gp7k2x
J/xFn86MgPu8Cvqv3OhxvLzL0teqP/E2suBoiODEQ/Q4vTMwyoj/eFOFFK5FrDXa
gYtNwtOugikBJZ5S3GPaseA/l3JfD48rlCxQZR6B+0Z2JWyI4OIn0i+Gl+k8u4vH
RmpWyT8Rub7iYl+xsCw+8Cy2L2UTLpV0B/hsGOJXIWyCbXl4IUNcQ5kEP2baUWsy
SwwZ5lRxulqrhjks9yaQBTrnE8UobEKuwGkZ4vVuIxmmCFMTTbSysS3ZLmBfFc4E
3jTTPQy4uyG3rMD9PLgjn6cTVf7/L+z9M6+v8+bsnJoKgwtwJWpBmBPFah14QLTf
tDio19aq7KGYLv0jnLquqkJttHRDDxnEsHfKP6Bjf/TH3BF3Ua/Q3lF3XLnLAYfb
zNnatk624HAyjG+SojNA0regkcuoWW2JjAU7BsyK1cRlTdckpvPGKRftzKmzBlqn
Abvsfz67BdvTaPVS8l/kP4b/G+Hob1EtlG7OGZNra7ZNMfMMkSZnK0u0tz6g8hDB
ZrN43PvZRgYmDsuaRUOZEY84XWjLHLZhrydzFaTKIpNNfwesnfV9lu9whR/JfKuA
X0H3PRfDmL3BmBiLp0+3JFPollexwiEBAZtCKTgp09LbXJYChs5bypMZMWKLQ4UZ
clFdKrRXeOGbghCL6w9WpUT2JgIFs81fo5Snw4tZwEKxASsgQ1whXV4l2gP8iGx4
9tMmf1vb2XUrJ8nXFgBr5JWIa5suxP/ANHh7IbMhzvMp+tlM9JxaYuJpkZu9Z9Nm
Kkvln9yqQTCoAHD+aJx4bRDFMDcodEDXs5czhPQu9VmdSBBtgtDcdJSby11kHqXa
eSLDygsSBJYcocULvItwnxyQ1xZRCnIfusp51tIMpwjAfsRTwePjM9UV2HaDMyi8
Y+ykRW9Uf83dux7lI97hSChIcMU9wIaqj7TvvFcEX3jmEueY1j5WugaqgCqNDBJ7
eWulgrp06XsyZeix7sSDxQ3JAwDvu2XYCQnQyZSBrT4GK6ciatzFoObCmLhY906n
k2a6/bFCZ5nltXRh9O/5hk1QyIVrmTcgm97Pw7TlUWgsZecfdi2JobPDV95GbzmP
HN5eAAVvsnBknqvVRb0WythmwLTUGMr9AqTh7opQRKi7ybwV+EAUqXolod9vPKsw
g6W09mQP3uaASmOP20iiqQnD5gBfO+c3Di9g3FUE6qfX5hjIUUDAFCGUiHGxlwq0
v7VtiK5eMHs7bzPIWH5fOiyYmP3HRiDJ6bRqMzoIDb2Ct+qEqPqaYYW7w7MGjrNx
FMPmxTvCZQYyZZl6QFyMLy/T0p9ij7OtawbueNhndWxd4rL6V0/hNC2SvI1OCRZ0
0aXxTclAJ0hTA5GkkDRpn+ezpYyQCw4VQngBW9MbhXm1bZYnxGid1zCz+Rm8ON4b
E0KbfiIXRrlu7WhWZD/64BbeggAFsAXbCCTS5kJubDlnA2ga7z/bQgunenhn9oaW
LUOmxzSP4LB+eh2gKfV1mGengzXiyYcOUTI9cQbkf5d61sPbC7eIH5z66xzIFydD
7XMTm0OzJthkl2AikaMPv3P+2/ssAindv68Gm0J+Vn3miRXGACipDNODNNjO3Pf7
WNXIMuV8UXlHvaIMlKIvSvtH31+MnI6tDt6x8y3Kl9y7IcMTNhHdwSsCVgYlNfo3
gukLmWIezt34SKaVoJFsqlkCxT9buk1l2XkW49MBSD7QGWAYH8uxc131bgqyOwdE
ThX3/ivlG0FSbjq01ffcOCo2T654gL8Fxx6NlZ+HKG2y08WWh6IqI/XRhtVCH4tv
lWcW4eN9i/Sz21swb3OLwJAbC4W2VExOLBpEEYigOEJYaDEHAVbQtg14FiGvFr21
RMN61PR32CyYmOgCeHSsXVfvCupFDuztT3fL+k51yOpS/l8jjqJzdIOj09v5/EiM
D9gt94KyCPRPc6amNXzI4ow7phVnYY6HQ+fIAN7P10ZPxmCzmGYE1clGCOAnWZje
GEO4Y9QH3cnX7n4/MKXxsDld03JagKKv2Gwb6AzRQx03jRp6lxff6j1Vklqv/jyp
LUGuRIieWKYiENCoSlku23tgKAw7y+eAum0ITi8bEnld3D3NmyjEvg5xWM3wtm9h
LJQxh6zDIJpWrNclIn3mWIl1nT3wAvLujXz6LvgtHZu8UEk2vrOLhNpQflA+9AaY
zGyVx8eRe1e2UZnPRTjrylsN6L3tfOuotyXoyvkFTC/lXfhIO7mTH62tKHpfLajK
Q2iR94WZlutupTUwdrYkuDrTdCGft+zvDJ9ily47T7smzMgTBWiIZE5l8vynn9Aj
aRR9oVhQP2eYAJUmU21n1IK0iMfAi7j2qV14Wpds07r/LXceKtiNz9ypXfze8zr5
bpqfHaLdzKYQJv6rw8E115Nnd0qJqdWfvkOYuQOkRhYnXA9B6LzluafOno5OIIQ4
DhzXN7S/t4ItiYbYEm0AqcQFsNPrV4AuLvV7gVgIPXnJpLqIaGymW78m50T/4W1C
trVErNLrHOOzhWLvrG9q/oLQmmjBxQuk8ojFljEOLdou8db54b6RumQ8Ji+iuK2T
ZsITeWRKC89x1TlbTdXe4PWVe0P3SrbgGVtQKMFJmy2H8LNXbfANjbmIVC8sZyOG
8v9k/96we2GpjbuvaLUA8K25BKlyyTQpZ7hCOaJ7PDI+FoAFCAoR62+kASqez2qm
0FFi0kxY0P3RySSCDQZ1x5fr8VDzW6I8V49vCSW2mOXGF2rDysIEdo3bTfleAs7A
nptS7ywgokJDY87PnqaSI47LLFPO5nECaSml+0VVakCV91BQo5Pf2wPq1zWNGUZp
/J4EbsDKojR4Hqxq0vOsgNlcw99eWdLFikFJIBM108xlobFgd0dltmWNIkxh6u3J
s+TP4UUz19peeS90usrWJPPhHK/dnABeFp0C5Ty2mhrFsBAgQVI6cR5k1QQXIVnF
oB0rdyaLyg+eHYbmpafBFQZXODvKWq8ADxMHJQl5ZXlvdsHRnKFtbduz2mrYaaQD
6GwJuKI1WR29KrlGjyIdArDriaoXRHZPxmCxZmZQfwE8Sn9NAUgy8fff6aDW6/LI
Iqs9yJOPfnduFVD7o2wsPD5Ub27ZXr3wgqs4LKwqB3SmKR7L+g5heC/1+JTbKq5v
JekdrNQ3TtMK113WDnq3wila/1Sp5Reiv6uioU/pi6YUyiA5BCTbtXTNRmDWg3nJ
6EkjuP53bHWziDgqMnwbZAb08bhWWi6JqVs3t0OqUUphtuJvwlaObKYIl+uF5UGA
Kc8/VmoiHuHqwlreVvzMk9wbV881EBv/BOmh9OzFjImDFyUhSEapFufQ/pBQrYt3
DRAtoad6EnhGFTIw43oQx8DS98V9ee/DjxUEZ8KADuDmHCjCzCp/fxzfBg5a9EHs
vQjKc7/DNlYK+MYg7avVSZuG9fWsmUzf5MnSMfcvpofvmmtjXYiptDnDpn6bpASd
1nUPTNmXgQ9jeJBIKaCFZfv1UJZx5L/zqVDVvIr+F2qv3y/u95z+NTTY7HQSN37i
+BHC2jE1E/rQE3Px5zi24BsDGGRUXL11vll1NH/CftoJbiBPhc+vU3Mkz9p9Q0M1
n3PLabPEng68I30HAEKSABpY1toHScuUX+K88Uy6wkNEYGOg/2LEHG66M/Jfu9aA
piFUHp/5MiO85Z/lDcuINUNkGuKoRfbImAu28QblrPmfcAX69qa59I9FVz06A3jy
O11D3txZ1Yr6AZnB+J0Eo0t/bQK6hvR/6rPU1cN/ykTg2/d8vdXEZHlfl+O2Ftwy
cOziBdczJ+wsaOaRijuFyroyfWpm8yZTjlZfKVgzByUdPFzn0h1dSkcxN9c3z/uD
hPLrYDFS+OE1num9VD94cAbakypfvUyhOMpxs7GWFykwsubYxuabUPzZk2RhZNnA
VIMFo4cVUx6JfkLVTI2Fq+/REBkrGA4Kz0j2DjreY87wpeXo75y5Sx8yiKdIUtg+
Irt3PqxC11eI1/2UdqTPU9BsBfOkqEZpUcBWK1lpa93rKJ2kU1rwMVxjojNV0VQ2
NjMSxPc+oMZG4G5ECX3MFw8P7I9M6J/icehRTxD54CgEoMWNYfYn7eg666VWFBM8
h4HIrWjCzyjC2wwLvI1bllJumPgxZPAVoDyeZequEQ7P8QVJwR67oODsFBrRuJyf
xC2LyK+K2RHDJfRNA17sswxexUF1qAd7SYZdsdViip5CZ27h8hRI3J5CDphU+bo2
uzy82VcoJ0QGMwrG8gjga7bPIu7RksAP3z91obmTYcFOXm/5QyOhFfIpK2isu0gM
LJfrRvyDkVcqU47FyFS95HMRjyApg5cx7v1tQMz8morKnNPREktZQMJrm81fJgA0
mr9ZDqmWog1LSasBGq6IJqyF1BEZxKjj7SfhPnjCguKgz1j9yQyntMQUOFCwaWDL
UEV8De2DOdSVmc4OMJdhg9rfTHE6wNpvbtiJj6EBbSeNjcau1xHFRje+YUkcOxGV
Kk8qUR2dneXtwp4KAZ3JhH+C0la15jMNGQFtixzC61Au5QWNKODBD2FVVuEszWRA
XVeG8ito/tZ7uFMgej56IPaiITabQA4h8sJ1lWbaS4JYx6T+y9ToyuNY6VxRHvS7
wACvAuHBDtISMqDUD8VA72rs8NLcL80DuBZ8CWRdoAWEpeF1tuJyMC18TAxfj57t
9FKCV/9l88IYTXyg5964GAbq58eHEZcue2F0fveq3CzjCmxFoC8wIsj4g2eR9vb1
9NGDIWhhnOC84Lm+UC9wF0KCu8tAGo5bjw9Y47WBarHfT7g5An3TelqqRG91hv7N
Cc0UX+DqhxvdHJZLMJrAnhdOtX2ckRTnGQyMO+ddpdmSzFC7O9qkx46qrqH/26ai
B9ySZLpfGYJLbXAv27+4IWudI68AUGq+XA5cPB4lAYfJRUSJAZJZ/JL1KOilKdeZ
X8ze+X4v5qeluBgXw1oopH32S2w3pCUmkwfxt2uCqt+3mgQVzJcX834Gc56ao5/w
1uNKqV0YKU7AMp/6+4A2ycA2BAoT9HAZUccaNGL+En39fOeM/AUpW+y9r9jLQ6mV
pazVxzMhYBT193N72rsDspk2p6Y2PzIU7+zy4Ce08rbPwNC6uQFbTZzWka91i/0E
i7+vlWtu5JNVStGdiGwFVZLz1PFA8NuHDaCaYwYbtSK3Rjkr9qvwUfM4GCRSqZlD
42grDLddGpaHJVRUADHOvGDoAjvMcz7+00QkI2LMHUFiu1f+jYi2vH1OQS34IQUs
jum+x6sur/Hfdh8NIuTc7e2iyZ4tl09s93DQecXfNxlLRvZGhXniUir0pgqGTOzE
vYB9/mN+7ENZA/1/gcf6gtmDYRJ7IzJH4xjRvYlUbqMjJrZ11InWcL4Cs9w56o0o
/vjuLl4D+fVkFxqypi4lKoF1I+Ip0wrMywYKtaKjKgM7grvjhVETm6S1wbNrjQva
nozYfo9y/uh+lK/WeUdKuZ6wHi+Lw5rLIoxCx8iPqtF5P2o2tn/3yaMHbiXaUC4S
P13MmGeDb7sxus2KHVsfA2fgJxvcpBGO2kELNV3eOjtYzdjMJdqnrRJW6aiqtrGD
wje7ap57A4sHn5sxBSOgitdRchx68nKGR62Cr3Npf/Pmv2oqXI4xWcthdqV/w0qE
TK5PphVcUTD+8iWi3IbCsRhyt8lBxh0DsJehnQY2d8vDy0jVbnwWU04Ck55t80TO
77tR3R8/f8v6Tr43nUDMRd4G+wDJopFIgEizffHFRsANq5Y6BmE4crGEgBv9ih6q
pYjBzTkAsZ2imD5DvOPfflm/FlzZrjTwtpXcPGz/BGSD+tDaU02aIBzgJwi3BMJ7
N0vsBXI6ph8B41ZAv/qum88iNpH77olYKjBemv5qhzBzV3ACcY5K4tKPAbDsZI2A
D2X07dwuUQ5ngnBCQR8FLilfRfyV72ViczsjYcC5R4EoYV0BYiuWjqy3nh34SKI+
akz5Qx14yRbWsVYtJ4JgVIORtpwatiEVFZcVwL2O/Eb68opNMn8Jgrx6HJVma4c4
YK1o8NwCCYpJKdp5S1Cd8rBU9UN+xRlxUOPIGU/lKh2msrRjP6yjBpJLmSoS2dY6
CUvkLpzjiq5ezWZ/EtgqTPBaJ0KW/0wbMYxqD5Rnd9rNO2IXYJV3ds1Ho0YJGfIX
al+CLyNpn71UqdrIXgWJVbc5ccA+UdYfKxilbUaMMZyL7vcUq//Y1YUQLeHjFpNN
Lce57P5knAqhaj3w7lzeBM3CKgqd8//idVMUHTxpWEKDYJm0JqXhg7GaMMXI3yvQ
QwZevG38frgnvUnljUKqyM+WLoBHb/nf2xbKDZSCo5gJ48v6MV1Y9pzvZQv4jw60
3Yhr0JP7qME2XSSoCQVOxjzfQjQcgDEu6Htg3YEmxSHJGzhxXyBSgv+KfOsEaQC9
ZW4gew8/YBylBIcQWMynNn2Mrp9iIMSTTmSlJqgcbmMQ+03+hIEmM3UecikUS1cV
fNZR/OOU167p0Uqhzus53A00mgQXhclduN2ujKiudU70l4PdVgRSc12BxUXZvdP/
WhQra6JSWj2WM3WkAX/0cT5XXRQULHhq9TTzIqapbKHRWx78hUjnue4X/fMeEcQe
+5UCuwIIqJ0dAGKLJiGEfOM6zotY7qLjXwr2LoXxkVnd2sFVtivn3dAvxelz5get
N7xjeAnKoMuXXZmgxrdOFUYbmBI9J9pbMSoussohcdo/TKw7uZiQQgSrZyLaMtst
bdOUYliU6/alxwy+J/hIr3HLluf3YpzEq8eFAPjNUJ5Gh/Yt/V92bpksvLRUfjm6
Q8AswBeQusDwvyfM7t8WtNs54DRNB9AUkNt1SN//MMEt/VBnFffcmSfE8oJojFIy
ayecdN3Jq/RenhRO3hNo8DvX4FBp0tVNPhbp2hcL6ggW6TT2tvFsnXhiNkinC+wJ
wYhfp+BaOlWegvphGZdhkItbj8ru63tfWB4QC987PEEE/55PtpeqYZgqI5fwori7
VpPwOYDDRgDs5jI2qDwCmlnUR4G86CXewmUQGyxGwg/203FoiHRbdnC6j0GOr/GQ
BjrSmtXMp+krxU+bFlI+wO0d11y6OUeGy7o3RGZasRvJ8I9Om6acpjtBJtVmlobt
eOqN9vl8MjAdDfoKmJC1hvPWRW+xiBvXDYL3fMNAJveTdxT6mNlP/FUbKp8Ht6VG
Fb5t/HyHGKCuDsbhSuw30Xepo9206fDb6nNwpf2bBZk1ve3yUbLkBT4jshyibBLt
80bKb/aUqTV3yL2NPm9MHlujzRwH7fQO9lMnqhrzJ4CgnQaRgNukhQnl7KgcSgCo
w3B3Ttc/yGl522W/WgPinLlI+GK1Pww6hkS6PQ7xzw61fweHYe/dovlh99l6cyB5
3qdrXjg3Ri87J0K4mtUZ25rGZqKpgLg7QObGla3UYtfENbKvcgtH6UUL1cxSAVT2
sc4FAu4ZkntdRhnQnpspMR1xZqRLA2pkMgmwKnBkAAqHUXf1tbCR9I/uJPYJO4DG
8qFhOKPIsoXzQGCenuUxmtdCbe+FGp5KdW3DoGHNcfya9vBlnhHvp6w48/dLswQF
IKlWvqpxXgzxr/kQo+ytYEJnjZVsICfjWA4CPc3yCrP/xoJqxCx0MHxiHvBkIQfN
jxem7cUFcNn0ercwnuAN3NEUI+B+m/mHMisxGmqUSFsg3rzF5XYBspunRfr7G6k7
5j7QKWBKRuwOAW58+EFRK4X/QhCWAOfEhvaCciqzLJo4J0t6qjhfFUJ0d+THD8Aq
uObLAazegM0Bbww+vrU6EO/tUhvGTor68MBDNYaWAFFadewn8nuFmtRKvPi44c5p
OPIKqqijfN8Xha9ovg+ffJKQRpWz5WIFAZ6fAiKpd9t2+HXlr1fRNSnMftwHVv2H
87LFNUtms6iA+tT4VB+K9ZjZx49Oh0jEo01OVD0/o6413tANAA32HgSeUN6PpF/m
jhbSR1PUu3ReUv28zZrhjvagjt0ZEDBudIpthayBpDhnKk/Pfi42HY0cW9Y48ziJ
oQSY81VgngNW5FKlrm55Dkfc4JGvh18xqGPHl46/XJevulRHkp59MC+4Wvynp4lB
Kxb3PtEHZc2NY9elYq9jOzKq7SE8gPzahXI4uCJ8C3ToXlOn7t8bojiprMG/u6nj
TW+d/PE9/8v6fzduQIH9wwrmKd4QQBDA+WWTM64GRzV73KGdGxv6MNy2syZtmWT/
ebFW6Oc0b8Rtck6vj0+aOFAdhk9UfaaRuhhM6UP4+TH/vO2jfeYqS0Yra1JvTlIA
M4qKclWnHzRosI3d5b0gwXXfJ1SaPWW26HerBXErsSuyt4ZqqzFG9nRsXrJuNmpo
f6U62Sy4FCanXTyd09MpueqhjQNrjWq9emo5cAxJS04FlwchOERDh0EOXAy5S3QF
T5Y1F1iWZlEpDqJeEfj8oq1NFjdxg31dCT9Yzw8hfVDhCo7lI5/XmeDaW4XFGEu8
Gsbr7BNWEX1Jh24B4dSGch/ur4kiQXDWR/oR6vTeRufh4qq9jcqWmyYirY6vcEhH
NQwet+uu2ObUSCkUExCuOjQ9codpqfaV8x1l+fPCJQ9Z9JQDAe1IGsL7GMHBIVEj
XKtrOs8GT6XdflmweaXeMwFX6eI/+2Xz2dlC1D66DWnKmhLa1KJjjVnAxiYVb9mm
WuNNPihNJjdfu6IURSU/S9A6A2qsjjTevOb5viHr0WPk9RtExbn9Y6atRN12ZGj8
EdpmnHDex4wG5vNt0XGEAbp74C5EbjUur19jqLTEiSMG+FHnHGIpLI3Lro6+nkKp
ZmsYfEiF8kSleKJxiGtM9wUrxzRUsIYivpTSZS7UxK8G/1C5RWc+qYLW2fn4Lthl
D0+8Y4A13H7kUsTZ42B8zZKzLj3eMeh7wzEQe1vRoH+kZa94YR25lbtnHkeZCRif
BQdIYIGVqaT+6T1guhaaOvE+/LiTkBxkjIhyzqZJYAVMDMr58No7Plpzddw7naqf
X3Qclp71JJr9Mmr5gz+z63A09B1+Fh4XATZtS6923f6YgeG+Goah3OvPgaQT5luZ
Udc6Tdj5OtwPn0mmA9Vpbe+okYMU0p9gg2+rO7YW/fKwaFogKZu3ncoF8n7EWCIk
oyq02FTKVOPnL8/tL2toyHQJKap2R53NLdQR1TIXcFwlOMPqwLrI19BsExZ5KSBy
Lx3SBFZbKjaPZljboLu2LGw0HxUIAQEERmoKPJ0LubbHzj4WDHD3SEHi7+jDNrej
hUBKcJeP6PdMaw2R5Uqn7m/4CvuUOtvz8G3ujIFIR4pnIDvTI6aKqLoHvNX+MkzG
SukOmrrK9Iz0y1WPN5bBuMOEKKz3iiWAem2EF8bcE/49Ng35tvPTbwyIuNulfRbm
SLouzxwFU+1Dq/R+uNu9gTYcXhmzY090kG/vNd5L8ZylVCkf+CPfqXUj2u0JKt70
+8m/swX80gaT4dVr2DoV6HKk2v4tgp5VdxWslI4h9Zcekf+ALZIFq+GkV7ftZaka
ra6VVlhGZ8gSQO95C+PoeIxh01uUvMVoBCK6PHlDUSyJpQxRKFOw/uKl2CY8S4/F
X4K/Fjvf35NXOFa8qmFem+G3pql6D9j/LTRnXHoT7EbS017VzeCwUFTtmAdKfjnf
qXoP3Qz5BxdwzIZZrCfJw2r+iDKYgYMRmMxkLLgNjZWKK5dEGj7op+NeKKvVDJea
Cu1LXIgwDjrIOmA1Ad/0tcyRuJQnGMcGCUh6YfsaIWr3orEl97Fb2SdM10N1Bglw
ND00ZwyG1xyeYSr8XpB439PgPiLxUMcggh/JtdR+/EVebk/0egKT566kxx5LBucC
RA7P1Z/EAQctb0RsUEhLTTpcAQ6cB6QuVBWL8eii0IHm7RBt9O6MVp9Y08AVA9z2
dY07d20pTHJ96ZQCTXMddlOnPi4M2e2qCTi9FbedNmTTjMdk41lbZAXN+3jXXBLS
xumzpcMDebcq6PLSyYmyLcCaVzB1AS380qDLOl3YfwYSNhInmuQzuoIZEUpqJlzX
eMtwzHwluvJF1/ko01l8UG5rl55G71ah281rk68yTZCxty+a3Q5znROvuTJbtqmZ
a2W2kaovq0fDvVRxd2nMxG6Op8TQ4gTBUsHTJXXVaa7/Fl9m6rhA/FMcQO5KIubw
Csd2Kf5Fc3P6YIIylNsPxwYQBsS1clPlIbzRKCrdh6PqyDU4bz6w/XDwNMYnjxTq
5rEU5JPcUCtyDFs49ZSiBMn24FcB2tsC0N/xIXXrwMm92IoBKevp2j974FF08Mw0
WRrL+bDNl6tlOPIxOWOKQvEDjHa3JV7Yws8N0BjOnkIo8uDxx3QXBlcQFDonppp+
aco/MEMtg/4BFmGKCFDqX5vE2q0qNL9898xzrQ/w/JNpm+pbsl6BD+enx/eSdbLh
7lLMFclkAuUVxJpUZaacUP356p9sFMLzqeGmeo/zBmsJ3TNva99dbYFbXnoYXa7k
8zWOHGwyDyY4VQSs4M0OduQ4OEwLaBvkydgjhsj2yXcbcZBisTbltZ5cFedFd1Jp
WM2NHyFDhh21mO75a66SbBOND0neKn8qvbAG55JcvRLxNXq8Tf+X7LMc5Z1rMV0C
PrWQArPkeAyRDUOwaJimgqu54agH3IyOr83WLm0r0tMVxKsf5JO6iU3y1yuyqj1n
j/FMYP41f5iwGPOflUxEIk8lcYBB4fCL7B/Go9xnNBxLrAj93soOlxZQXchRslr5
UdB/96d98kQJIdES72ScuaDcM6eKDDjI4+bIlL5Fp/KUBCD/BUEcOqH+qBiqfePH
IfE8HLpqyjNn3x4qAXoYcMTyRkZZnVyM73XOYCtI3Da6Us+fScN4X2vhWzWxA3Cn
HrijGZSMGOv75s8CPPXRupIltq+9b9jzuZ/0+YT69XmFusPvbZFh3GfAcngBCVGM
bn+zGZdE6JvVANYPcT0SuIS5v1zaafpT2Gdlas6vGo9KIcG4i0kn7ArEzsHJUAlX
C6dLaqd8P9weMjPPcKZAz7sWUHUlaEtGH4OqlpZ9fyrkJZ83YuAsAekNEWnzeHJD
Ye2I68ImKk0e7zLvp6UBCw4r58v4HGmCjeq8pGJ1BP7xx3VoOhHHRCjqCa+Ie2QW
RLlmQILWSnl6IeCJgGwqIHyhmwSL5BxjC1i+kYdF6G3/101sWWNpd8FElIBpa9Ee
QBUSuty1S3Fer5GTuhzX9kIIY3X6Nr+alBN5hjQi8JIRq/U8AqjY3nCOWvtGfkCC
5fBlyCL3E7BGdzBDUSXcNR/756/M9p7m+Xq1iK82HTQLF26z2j3jvw5SF+EsF8iz
Y0LdboDKEdy0bBzOl2Za60R4MJ4CpY93ofsg5zAV9j1KQxIKJIbTWj5yAcSSr02c
znhmP/SNRQbMWIWkAnVhx6D5iOfFLT4+cOuvlcs+rzciup6SO4MnHu/Le7cLm0Jh
DK8YaGeTHso4pPdIBK14gNGqmqHSDmPgXmBHRxNGu3KSW4OcCVRi0hkg/AzDyvFi
qQB+d/X0EOWIT3fQbN35l/wRU8FQY+K/sxaQwrG3lRKqjLrtyU7lWFh3+fnwKoo2
xVzVEQpqUMm9S8ql9K3mVARJGXWDvzcFjVt+dxkjkZFNk8W+9NRRwNTj7QVdFdaw
0DI1ASHPlh9mPS/HcxUDrqEqWELOeq/1Uwpiw2faalgKvh7U06Re+449WH1KtFCV
OWDRWzxKep9/zAJCfhC6w5zKGBwFzkYuUj+vKUyRMiTQHemi0vuFMxyZKqmKxqet
w8Xzr18d/xjYhfZbunkf9IsmH5Pf62GR8r4pKK62uQU5ZYUDouJIP/2l/9udHKFc
oe/DPLHGHRdyK/h03omMvQZDRW4psC9Q4CSVP7RhPPVGPOfyRaEtMAoakwy+xA/t
iz873jG6hh9Eplb3dJL4ciGFXYpp93jEhw3RIJIWOFaHclivZG4RB7CydmUKJ6jH
W8wuTobJ4xu4HgxR156VVCIlV27Ej6bx5pICc3sjkMVc4UbyC22VREAWIR2bPnCY
kNVRZZ4Tpx+pWF/LepO5FU33AtgE76xBp7EqgCq8NwA/JEgC9smqacoqBFr0Yr6s
MthuyItbQdxbIEuP2Wt9BoOKfMLS3nyarBJYyIr6GG3Q1ZPPAmK7R9b/DFPfATqE
hbRbqFLlGxIZlgEyNdhMjlf3KkkmbEiAg438x9pl6iDnLC18CVWrI2ZoINzMuGOK
3440dtUth8wQWZ9U0eOUneF2RC/8Z3h8iXFhOBSdYyEKL7J708hzu2kDJyCliFOA
QPrEnwV0NqdM0ghpk0n3aqvF0fBAUIYRwAVIb7QQ1UMxilFATRI6SQLGt1urL9GJ
Xd5K9YsMUjOaNKWJ3iPrmoE3S1h4mDV4O3Ahyew+shBz8FFq/mpPr25yykMBBJDB
bBnIbP8z73F3JiJ2h6xKCmYr0V0nXR1DruVk5BtEfKtgn65oxBKpGHLU1r6v8BEl
0WVtvb68mqWG6F6IPbc8izQ3g90omLjD8fk+X/HCIwAZ2/kp7ZR3EeLI/DHvlQBH
MhQ2lz9WTXQhUiTDzaqceUyaNmaPyY4uTk4mzZWSM/gkeePjubNjka5sdSrrXKHW
BsIUzpdZwT7STMORcqmAhAifrQF+SlMF5b50TcfqSmyX7KcdQOLop1OLIvR7KHYb
07as8+FaMrHoK6HqNk1DqS8VQCU0b9kGS5zhG9obTexgK/U/5Wrs3EqRIRaBBqbn
xVUt+VKwWPMWK7s7hWLJiVSUKkbm/wqKt8O3qLIWaHb+iAzRjZlrfz7V8QBvQ2Zk
uT+a1fmZo2YlEO6URAfCHSmqe4Kb7ne+Y5urUauckE2IWu4EtCp7pK8AHfJ7ig67
+svU15krWS2roBAUMVtmLxN9iSKuolDF0/W41ivtAXUHX/IqoApQqFTTRZWCePTn
ZEiPv8vi7H8NjAnC71BKItRJiQLbiCdzyNdG2S44NTQZxV6zCs/ER8+Sc5Yt63iW
8154VvcWd+SeU38sUlSsU2baMvIvwiqfacGy2N8nbdJnZz90AR0Le18e7u9F0vlG
LlHTSOV7NIQdi7fLXAw+AU6nDWKObh1kGeOWkP3yGpz8rvrMQ4vWzf+LqNzYG4Wf
8o8jaBqvktcCxIpxJHFU6QjDo7TvMWMTGSecHh64Ts90upLVxm4VPm7fWT55oC28
ijk+H7FHCA+tieeqmG/4rVg7X6Q7X4dGO8jNwCyJ1h4J8UMlR/1qOfzedKMMnido
oXmVehfBz3+LYwBgIu1UjSEKOg2b/v3sExvQ2TxxM6Mm1W6SE4lwVpqECgp8INMu
kJa7qr5OgaQ5zSTCRCbZO6hEV6NU8VduPrf8odjiTRZZnmXfE/WqwvkKxt/cdMBl
cBPWDmoL9J///Pa6ASCsK1iD+cIrqZxEg52rk1B0PKhD4ABDbQ4kH2oyv980g0jf
uP5tu78PjrDl8t/0KGrM/xHrluTLeE5yTFV2D5l7UlAUG+xTNNg90nFPYmQSEa4w
TDCiwSUUqpXarQzXS8XmOvDquTO+ALxeaD+vFOHD4wCdgXEwELThYz+HXw4YU/Fi
nUAxTXa8RZrBfA+14MHPGBpJX3ctEzBsAWxHuC6fLoxuXblbTpsYchOWE78e3j6Z
aVYHxjY/0qvBJf+bK0oU4fQUTuAZt2vfxAjLCwvcpa7ed/bBixacIb3clcIQ+DGv
ffylFZoIP4blNz5CfeoKy48gZ/Dwv0ADgglevj9ynfUthbuNL3ToOO2xFfNN/liP
7SzGgRF9h+8W9br7d5Nu43pAcuCM9xQ+9KpMLu0gpI48FS2JOYDDy6s7D8RoqCBf
FIWQ+UfhjwezhRKvEibQVSiaycGLSnl3C+VQnecXX1cjKu+1247T9vD4IVIwuuft
tLI1r3BIxS7yNEmrYpjg9yRsGGEcjsWyNZ97q3rZH1YupXXRyPagFgtCivNA0keH
tq4Bd70BbU9CDOH2CZndUOUK9wbut/L6AOdDE6+jaMHW2ijBWJAdViju/HpUwmML
9/0lT2D5iWplpx7n6IwzVthRK0AwGAHxca0V4lQSP85e9iYivBrmbOX4Q/L+wbpk
oKsuom43e6OTOh1dVu9ervP1LBAhZs0kla/mdwSwBmDgVus8TFodOCudid+eKzZ8
tdcOnweajkvdnXwsbR9oNuMeccZTichhipK6urLZyjlATiNC7gg+B6rzfPNxDZ8y
dW8HudyAYPFG34xmPqNmaOrVgZpwRne9lC/rF9At2K3PfnyL0fXGy1FHuasmsCrX
ARpIK1mBFvGDFEQDgPxRRkXYR5jwyRt3clM24akZAGTZKaIl30KRDFDFo+BWfiRL
EioE26NKSZFY2IhyhNIFXD4gRsnyGZD443nKVBabWIBHvuO3/K3TTrsMlbLYlL2x
s1FIcpqJc3IqFTWEnsRO2Xp/wyA8XeCxgpEelNhwyHBzzvBzE2Y0SL4kalVhHRxN
NzBk/FPQsUn4hL/BlzlulpmClFVHLDeXsP1gQ6EzZtJlIdykbHsDrz5hNEOvD+a2
7/OfNCUPPpYe3tJ1Pr5H8TV9V36VTcRUuCGqe4agplrxR/xQmYCDgiw4GcJLG8AV
QlEvJoTqidgjrsZvBk/m6xDG+o33r0s4Y4s/95EyExxKbN+yjzMvGSYOmHkbPYvP
8pPR7IUeiosF0glE0V4hOqUQL+9vH05X95IoNCNM0mt5659MfLSR9DUYBk9+MFyQ
cAJYakllN8SSetfimkOuivF/Y82Q0iTcq6VCLvx3QfDq9jnNavq6OisBMJyu4Dyg
mwqeEgExWhm+YC8hj6hqxHI9d1reT43swuHoQI4K4f2FL00AP4c4YnHRJhJUpq3r
Aojt4iTrFOpZjH0xNYQyzZRgk/X0S+BpYn6ITyKwX5OEE8VewadSikOJfkv/sbGn
077pvWZe4Y/fwSGPSqi7C6y8m+2OR7HoEX9FaNiDaEsIHGMSjVZD93dRLt5Yl0T6
bIGtrTSXI6cHkLaqnYqon+RX7ykfDuJkABkHYp+6RqRhM2Y68CawNsxerhVET9M7
7KicCPv5NUAafxO+RrIQguS3UMmgZ+4qdgHklbed8mJ6LcB2XQUQ302L8omA0ldh
a8w9cUwzb6cqCWxYZic7t7UP5pj04n+6/C1+OQ138xBWXfPaDgA+SR3/sHyNcudW
k09r0VLvv8e2SkwB3+PMriTXQmDiR+u54U3erGZXlN12JSVN6ahQC8OYwdDynd7o
r4uN6ET7vY/693z+IPHoSq1I6Mg9rGgbLQmpW4ZKwDt+4NtPvlZbk0q183/5rCef
HZKtPAJIeevXXjK7ZNV+rEVwE/hn+Q0MBIoW1dNiGoav4LHjxk+mChvWx0rsyn7q
HFl4wyYbnq1hpKxkHBywcY4/avM+Cx322sJiBL4sXwjWvWdRc1eCvfOp3gGCVDZS
M263Oe+87fC6weQEg6hk8pVQNBJJC6qJqQmBZDxa6SO/PbVHcvcih/coAs42RWkf
/kwH7kaCPImWlRyiWCP28cut2w9t6d/Q/u4wxVVOLB2441kmExAEERqje0qbE6yv
6yhuLoFJge40PXGredBH8p+tvZQyUJ3uvDMl6aUq2lWtMMBNKD4nuqrG76727fXd
43RVgNc0mMj4R7ZgyTgwvL8/U8hUxxvywAUy3CeQQL9kUq7KLmay1hH9ezY02a/a
9VC66IINsGqX69kmx/UFhzfqwORCl+m3W/qIuRRfzZl3/aBKlft8unmqc5zJIDkT
K5dyNROSgTkA/9sSaHbcUOC+oXsl460SSCwGPVvxBebGy1ytik8jVxV2sD7DT2Zw
uxRiOVq05cZssBaU6FK0qZz5QOphZtcDgQx6lmMsusCuyUWIwtNSVYi0OhJpoWbz
hRMrnnNSgpB/dMiwtqMQ43JQecqJezlaXEGWOAjORzDrR8knjFwzFfeeavnJtzaf
6fF+xcfrS4Mz/IfupylT97p/2uMfH4GQq7QjG/C2l73tXafhDQCwmmKdNJ0f4IMV
ombmWpDdyEGUs4/6C1NUFY3RrGS+j5/JdO7WVhZGxZNNBwMaWx39gfxavg3nvcX0
D+VQFbo3dY9fya+g6BoP1Vj2dTeuh4hylkxurUl7zK+2Xn4nETatSmNkHwZBFa53
I1RLqfqerOSNlMBrrxvrcDubJOTP/y+rG4Wdt9yBNz8ciVcevjyfknkKmieoPY4P
QWsGqRdyjDVlFbBoBSyKTKXmM6WQVcDlBFWaBUbazSTGm9qYD0eXjHdG68+Dxzov
6SQw3BzOq9AY+WHF0rR2EolxABMb5GSOAlFnwuRAhCWdcqXhENVQauwpg3w808gX
wywSUVqeiqNORF69eYI4pDUqW0XYWBytea+LdFIsrEcYh8YOJg9B/E45vlUqSnFH
010n3whj0CXM2HOWC95akJSMQMKJXrKDyHiHeELeEv5S2pI+AZHXrvJFeFpIFt4Z
sFXqDbnd/i+tQCQ78cxxNIZ2yjZ8QXjT6EExIEPob023Yo/naIWaV7NPOw5HK8iu
voHYFfoqCPjNYwVe83BBgv/qOVssORG8RgovsTTwjIcROQjmK4hlLgcyXZ9/y6xK
Gq5+6ryHsmmf09+ZBQXPAtQzs9IGBsTlw0y8ttRM2iPvlva86JoQZ1Wc+VXBi9sl
QpX9DvaXLOXh88kS9ODPB5AMAf0iA2BDet3hpMHWhtdgnXBNM6AW3kfRsSxv1RRv
ruA7WOtq0xSdWvSRw8ptDW3I29tnKzRd3zzhjLC+jnx/MX2brJYmcJY+zmbDy787
hAmoWyeqVG2QOLfpx9CD2JIzAEiBOR1YRucGqa15W2XEgTVPpVaCnWY3vVHdUI1W
4PE7mfuB18UYjr+MkXMCKNM5Kp3AKbj42etatFHi+IrUu3dBbBiHCzUolVWVOzaC
a1R25hZ2FJNGh2y6c3x+y9lPW2ngf0EZLdotiW2o53lOmi1Et+CmPPorCjQCRstO
yBrvXB+OPtwash1xtknEJjLJTvhEVfEqdkcv8wTV13yy0V8i4feOm6YsC/KEGpTv
kbPJvbz5i4/1yiLIYMu2ttpTrXo+dR475RXQe76W+s9hKs25AkLFQ20UrGwZ8cct
8J/02QlXdD4SaNqaQM5D2Nbeen1A9Y73SZpyf+//oYAy3gNrCzbBs7bYQ+cHHVi5
+IMmi6MUZIwvGbOrVu2zBy+Hk7ftCAEPRP9VbikL8iP0IX2nwywNGw35qJIsDVqz
5ZBI9r3iBH+TKrREqpbnh6EO9i43lRcIXT38vCem5oe5NqF6KK0oSrdMbDUyLjwP
LaE1XmSu/H0B8MzwFUlCePKdQLrcz6bL18tzsYEPI8ow0zfD8Hx2zow0c03Fk4Wb
GPKm+oIVc0Trl6dDfg1SOTNneEqH9zzUr6aCALUorgcGKjPxEt2QTlfKHNf47JyF
Zy13ZkM7NrqvuiSlfTnOzFbFsmo1AwlbBdFP/4Gi53LdGj3pcQei4ls6P5iywlYd
5gpMSci9UJyJktPvkk2N6JSoxBGAZYyBsyS49XefJWRVXaJkFGMDGxhWmAnhTdr3
P2afwho6r1iqhaHAoqS0JHDQKyKsaJnDAvsSVLv3Z3wBqXKMOe/PjSngpAdUu+Kt
FFCwDBHNPVHYhRrL+GPcfSgVTsGUO9WFh2rbPVFoGPtwKLY5eu3LWTlH83TK5Fm9
w++QL4Lt9ouii9Upm+RKrDrXsJYvotpAcfr4HrpcOHTmAOFxGeuSymESLZo/vT5V
3jhJTHEnckavhSms3sx9Drs6dYyZvIzeId/tlyNJF8k34IWno2F1lUyt1RjJPq5+
gtlmXF1uHwdLsb9QH1JNLD4zbSuZKoR0CzXUzEm8655FKnrxbBaRu5lKKPyK3rTb
UhOLtc1f2Pjs06uUzSEjJTio7EZe60EMIULhNmT++AO72IKKKzfwH6SXYpYE2ufO
MdB8MOzo5Ae/s1Y4/vBkxXIav62xQISo4+kdwTd9wR6tOWcLFWu95eYPQUis4lsY
h/K5bMGJ/46JLWfvkhWekvO/gfyHTBZmzFdxJ7t45sQClXlRX3NoZhkVWVsEh57o
JTqA1sMQFtbQAHN22qWJiqsP5wRTp3EF6dkCS+6a557tnEKKGlu5jguDN1juX6E+
YSElMyCa/W+Ztr83oiSNhZmEO3o4bvnOIc+ZmgUm6FLgrkmD/65GhIo2BKGOCoOj
zmUIBJ3hTz1ApOMwihZMaMvhh0j2X+FBFKOSpRbML8Dx5eikLY26NNSPb0b+BHlW
gTdlX0h6RVGNHvAYzTnTYW+833XkFlP8qOWA1zXS4dbjcelJgPusJdMotOqTUk6Y
ORSuHWtF8KpPdQlLBQ4Rp+PwLLy9BjBPitG+cu1Hg8JQrmba6O86eQiKxfyM6GEK
xCGGI0af+wEulxKFPJe2gRzpHhmCf3bS6M0wBPMd6QmOnesXlSqs5bOetaVpoaR5
1vZlamHJimM8TbRAdg7/HPvwFosJNmRJkI78yVQlxUMG+lQ6pEK5+BYf41W4yVfY
bFoW/sNATO2ATVv/yywFKNGmLLzcwiCB7QG3sqqYEL7SAD1uU64i3ggTm+Tt6v+o
3kjr0c0SFY8ux9w52MVkTIOpx7WyDZXktw8slmBNUn4WIdS3XQmwR7STL6py4/pV
+rhgTzTm1tbNGkLwlzznk77mbCJQ9WRE1tO+XiCDeqciXggxYqk1fEPjh0AA60kP
JC5E3TQec8Q01DUD6NRBzCOVMFKTpILJsVFr7ht1ytpLNGer9LFPz/dm8NGoje8T
xGoxhxVXnGtrwDVGipyOfupslFyunG8RWCKxOh7ecaBrWVYyanxMZqdSMXGlVJHa
n0NhFH6qZC963pb6aoqcD0QmzsLyloqElt5Ta6ZmP/EMbCKiv8nXiOpXE6h+2ss3
GxLZW2W/b8GQNdXiQDryUdJGqAdXDZdnc5S8YqxSOJvJuONHBib0c3fJOcThjkq8
RVyAz8/2NhagrdkQNgqc1kiA9C3f71Qwn10Lh9bjWqyYck1OcXXQBgzypr4vW+ca
2V1R3dnC3RgKKBY7ToNGAk5AwsY+2/tlsThkKwzKHmBkuOD5fVo8wnSE9q//B2sU
px+NeGn9r76+Ekm22bBMdEZBe0n3KqZ71XPqV56xYiCualzJrn+RevPpZka4l0uu
Ld74s7hj5+ryXkYmf4RiQ1v819tv7gHU3GZl8SR/3Y4ghXBo3TV8gHAVhGUsAeHn
Q050k/Hxb5lH39tG6TXu2k5bWkGHjWFimeZZOIJDSiETpJhmRTL7HQxj5+vlTk33
2FvxLY4E7fUz9X+P36Rg6t4aTvdZVFbWD8BKfZXJfqFh86sHPsPYuptEjUl0WTB9
cEuk7AUj7SQ/EGj3XjRq5laLVgT5YPWU3AuzVKqSl+m6m//pL/xbAzl08fkQuNCp
zw39/aPeCYL8g5656eGrD/c2R8HrFnxF9DWkErKkOyuaG3z/+DHun0cjfDBUeYko
XBVSyKokCzaFe9mfDH2QLSp3dxWgmnNqwgxJmfcw66XijnHSHC+/vCv4v5Zlx70i
fcif1QUAp1V1QKnHWfOlLOfAG3C5a55EFFiF0NPrxE8r/UAWDqXBGbbz0gtPYfbI
pmGNix6MZNlstAIDPv2LXecF8fsa2zFtdMO4lgLJkI8XNTGQ4gUh2j+u2Nu5xUmR
sWKmqkVUQgmgY16qgs3CHc/3sCGJ58FuKD5mmjVEIvK61xOxvuxMzrdqPM1vgVpD
Y8hf7pRKAsIDlq25dVyt3u0GpJYp/uj942O9cnY/gWGZNI4R0bmbADHdSEdQlqGl
k1U9Ixr5Spj+iTVcNDVJNR1Pk1Uz3GAgpr7VThxeNf8FnYFBhmJ0qOSH0g7PgzMR
8AF3gDvoyKBJ9yPHxRMJ78qV9KisuVp3JqS6emAHSi1QwK9Y8OvrbRutTgpzCA2d
sU8B0/p3zBkzOno4FvVDDz/u3JknLtDfENl3BNJB0C+hP9W+g7bKMnruDwWo+LSV
kqh7O2k3kdd5S8mQdxzs3uFcuBybfA1LhDbd2e96YxApgJ0rn3Ivjhvydmuq6HwJ
f2k9ozz6/Mr1Afw0H4J3ytvNLh4DccESjg+P865NjZMgKWdlfoYubEGbjMNLoACl
U/crtUpnQFgvAEbmBOeOyCvlOee1odmQ2GgWxDRnvNkcPUogyCptMU/vYGQjJuDi
gCwm3BHcO0NJ3dRxlXrZH2QduCzhxuUc/wLoiRSCL5Z0cdCi8RdQLbDVxDFh8vh3
AqER10dLzEREzwORWclTNHnfSPLC1amJwkvWxrAM0s3idRSuvMX32kaja8ybzg1x
GgzyxcZm/UhK7+tcHEDz0212jXH7zbc2njlJ1FLtyDVh/tKoOcSgTs5hF/12rC6U
6PNmuB9oJ8XbVBV/MEqgI3Z29KHO2c14GSzYEn9ltjhIY9vvdu7zmr0sJYcr/KjT
ENSeIRzG56HDdEQjKov1LOoc9mH+125Ds/KW4dQawk4GZEbZVzVDJlhszMDv5Re/
po7yVLLVlxOYUacfr7Foi7yneZl07/hP5lo2ujxD/b2HYLn8+ttVo7Ji2DtZkEd3
leqhAuF/HlgE+kSOs7rENZRC71g2RV1D1c4Im8KP73zHBHBURCaQcq6PjwS8InxR
iD/h/HIlqC2cFf7zgXVfZSnQhyCdyR0gNDMW1LgwcpbieVfZW5VGuxiEoKJUawMH
gWMjyKREBfgvZn6lrYOTTZtxbofSXt/Fmepcod8qt/Myb77jIM+C7P2pYCJEfStD
c9bqzGG8KsQgPruGu8TGHop2OoIOIclyHUnRDcrsP721MyrY4mITClMPInon9grl
p8SbWy0Ez4Q4S4OLSKn2OjghNpGfApeYv1d3P8N/xYUH/i0kh5xwVcpyBQgogfaO
qN08cQbNmFyhEdxkERdEfzFan8peaS9lITvE/SNLBFZaCency7z+ZvrQsxdStGGl
spEQvfnRz7TSumK7vmDQJpSTF0PpyAAMM0U8yhVqb9ks7EnJP/H0S2Ajz4LKESKa
mBXdzCj8sRgObGB2dTZx094eMolNBN6sz2pP9x7yBPQrgUmIKU7EiX9nzBOSj/hN
FUTd1o0yUFgfMygoZ2H9QRLl/P4giPfYGty3D989KPLGhxoXSMt6Hk/tqzRMBJep
hsueHh4UP+nO9QYd3/7mW5GUxgRdWj4qRGocMPT4vLVuyUs11XJGuHsuJKQDwTIf
80299Tpytz2GNHQvTOT+54dO0JThlrTKaRvr27zZJ0kPu/YOIG9Yc22W/rpR7KfZ
Ktxk2sr1j3wbRh2JzNvaJjLOHPnZBMwAUx7McLokMBRLumBukqF+ziKd6BEnoSV9
0WYkHqW0JJeArpd9+lBu6nIyV06lzzKykaGmbQUKKDtgUFPJhg6Vxi3aqS3UsAYn
4058VrhUPHNXU4DDudRjx1hCWY3j9egv0hUBanVTz/8a6tysVu7g596A0mMHKmZl
6PFBVryomC9JaPpmjOJecfdMH1n0oZLVkUbVOGDNwNptWXE1Rst6bubPoroY0TOl
RgLpisUen1wuEJEYKhuZBxnfjxuJbGUEVhY/K2KlgA9U+fNAtu5bm29mBiVWQ7Up
odxGvrfrtJESc2zJ2trcYzmpmsjFSJ8EKgNVJg4g1qeBAkN4jYFxUXznjqZVy8av
HcQdpTG644NVDpjNBj4pqwfApWROww/BkHyCrAiPXRq2GRgk5tFIo2Tt7LLUHE3c
emv5bxVDV82rT4ayuili9hVc1Ypu+zJ7ZqPKJTnrE/+HXwF+Hnpmo8Mx7okkZznr
vqrKv4lvo9yhzhYmSkTujgaftcUTuAQMLzp2PnOlRzm7+0vcddtp0GYSg4VLDU5F
MNihac1VIZ//7AYGojKZUSUn6pUATIdfr8W8CUWEkeXKP6BrXZrAbaMAR0jVnLqV
Ygs5u4MEuDW1qxaCOQCIn4EaTZQUsoQ3Vfb3mlsq9vFJtGhs/RJ47i1pH8AyH0kA
huTJc0QRXYB4BowsIqQEqEv7djBS5crophaxskiRhyDaUAgG1kETSYyO7twuFvLU
pBT+6ZbhKYDqvYeBy8S/aet/RnQWg9Xjx9YX8ueb0pn5ydcopnH/A5dVin7RYHio
iZ7gFLWIfiqb33sGvk5osOqJg7C8S8o9LUew4VgzfrVqtRLj9CHNdUBncy0R3pCH
ke5l0zxp+rASIdg3cBhZORIQeIcIe8qURI+ghoiKra0gBDjq/Vo9q8Rm3wwqsB7Z
8UHUUD5GF2eS0YOpoqAjwUZvbGMlQy9bQqG5YCYFghjEOqaU3wwuqfHU2vOlIZoN
VkYP4Fx0S6rYrPi11AcK370Yn1gmabBjnd4u4Vb80k/aD9mJ3itS/ooqHY2v1uMH
2ghBziYkGrofEVIqXkpxA8lflyNgKUu888LaXyu9iJo6KyqezAX2zxyQO9J526bE
oIh7aWuHR4PGBSo1r+sO8j7/llH/qt/xGOJemrPjMN6gWwHkKaum48wV8/yw0Tk/
ruOvGpxMBHmORinYsuXKNAw5EWzZi6plvIlMyVn2rGGeHlH/GivcWV1K4u0fBO+W
ACNLSthKPnrRUVKeZbL3HnJFDiZgNMmuLuZsXiEyeOPoSdFdZsauwXjwWuIAs4WM
V3TCXCIEQRKUlDZzRSjUKd6EkTe4fkGXNGq1brhVQS8LqSFghPtEIPfYDtPXj3uy
hu+laB4kG8VHKFg1L7l8Cvm2LGB28QOhMXkJ+z7PUSYnMdbmjwtjsqiWZ3L+fwTS
zwaonS8vmbDCgAMgnfRWJ6V2vv12vH2O0Mbmr7FfpjOpM4cQYEu5be2T9YJtQc84
jNPBVyeYeawSELWJMR4C8li0fzSTMbJ0qAON/YGMWDfDwImAoTFFF7IvI0kjxuGC
UC4rOQGWPl6WP/cCqHNOYaBy8+HQHoznDTQklM2BQ3RxNMfi7n7YDgE1GInF9fM7
vczhdIUTBhHO1UPHmBlj7Izq1/zlF+qF25jKTwgogW/jmVZSu1+KFkBR6lWKLwbB
ow1ovBtoHdKSdPpWLGMfi1MP53RTBlCF6rbbVlot3DS+rxSSAoKBdfDDsv13H0j6
Y32UWlFDVJRWARORgWPyac+M3O8T/haZV2yhBshmLJpbNmAH7isH7bAoD4UxinZ9
6cad0ulmfZBSlq8wDP/cU7am7oUfBGaU6bohBKzOkkq7DUwGuQeMGAg/Q4VC8LTZ
qrPyKIyfVGrEkiTpA9jFgk4rVlFm+QuMI8GGpQdBgUk1PN6Ji7BifOa/s1ae2QPp
9G8hNWQqqAGmPEw+Xs7yhP1Krh+0QGiy979lw/wbQ+gsS5WIjXxCgT3vqkUj5xDj
t2IPBq/AuBgaLaKB9DvmTCVeGvBhc9PmefF2kLPB19JPI3FMFnG658P/FFCQV1jw
L0Jzd42c8PSRavbcZaS9xx4BZG1PLs8bCDQP6Ak8aOw9Y+ubXyhZp5QkfeLXU3VC
Jwm1ATSK0OB1Y5qw163fDlqVYpR0RCpNL30cYPhs86mSNe0pTrprnaT7ptadCXQZ
WIrQcI1hRvrsXScRSlsSIr4ZGS5U98vLR2eWiFmvi+a7pYW6mRh/Xe87o52QA2TL
oVebpJJl++cEXIOSuYm26y/LhuCZ4oMT1zdFSDHJFab0jcNE3wbEj5QEica2yyF1
8WKq3+1irb+XjjGJ9qsMjZN2zIYv07rNPMfOzSKRU4xMkWUCYKl9vu0uFrtzbjVk
lwIEYarfujCsOQqcdgqeUahwszhaH0n0OmhR8pQep3hkUFKm66q7zJFTQDuQigyW
jJienxz8bgVql6uGnHOi/acsYG1rzuW7ppqV+npqHGBkZOFx/cZGKgyVyyKX+6lz
LWWIwKyZD9hSHBepkl7JscL1DdeVOMXdFBbMPEYk/6fgWvlTAy9W6UmyRq8xcd8L
IAYZtoDpzPgJqL2lQt5pMOHfr1vjcF5FbMTGVeamykZDr7ZC1IK0kBEMl5bAnvnV
HMBVOj7eBrikF+2TIjICwjaRDq2fVMAaj3akLzzRg4d/jYFrtgSVmFq4l1X7qVbD
D/tnNCsTq5Z9XzrtDAahKOvtaH9yUee+OmrhLmClfoa7Tr9/CU5esOMUj5D3wAil
HL4kAGa1Jt+ESWRX9zEEeLlajWV/ME6eOVIzXCcMS6vau+L0NoLxv04KxiB7w1fr
uODMy6Ca72FB23vQC/tSNqLbu0LpRixtFmBEkXkD1wr3IYO/oGegOryNX4LNurkq
5yaf+FUViYbdSgInwPYv4N6/DJ9cX3h2kVlbYRDRVLvYKbg9bNE8lFzsBU79e4DM
ZrhDTUz0MQHt8NLavyMEbqv45A2wZS/L/0qAMCQjZtyZFK0/vPIfl1KESDMoNSiL
CjrTAZXgdxBfNr4TPAzPPU+2tMGi9C3OurartffiNSLzVeMt3YooygacHZmZzZ7c
8x/yyFmLXpnwSv5c1UL+al6ZZFJsxoSV1KDEGVTDV1ziLKpunX0z81ucmIwsNysd
rCzQ0yd2QZMP25LMi8f5CHhhZtsJdbrlWvMIINIrzjkEGXUpi2bGE5D+/k5m2fSd
aHamU3Bhl3Shj5voljiUQKwhS6nXQVi2RcV+eZF6JiIJeRwwsMY9Cq4OAdVEm1b5
ryiyY4kLQF0tflAAl5YAzD//IBur2n+eg3Qj7Ozel5jEecpK7AC/tmzeUjTUIMd4
TAVbO4tznn5zG2Zpa4afgVo81A+HXiCIXhelR1mx8OdhL8wEtGeI9rx+FpBOudfD
Bh1z9gRQJlsTsllrKBdrg0gyVcW0pclcp7UtSEGdJnlk3ktd7jpEyyVsAcXL1jRf
6DeKTaD6Kz+7Q/NngMuur0QCYTfEtvP2fYmkvdorcKGs4Oz3lBXN1gVOpkk3vMKb
HDEPHlY4VeThkUTqgufxj8mbV7bvVnWbbsSQaKuIx9+rFLY6A/HbrHUOp48Btf4+
Gv6Xl1ipKFyTsdeRwwGtwbEsr6VY5T9OUAmhxNRrA1N3l/pcXiP1GHbxHm9/ZU3b
QeQcOoR6iEXqVgfZ4HOgpLD561Cvk+wLobGASn8gdy2O6CCv7UEW5oZwBqtH0d3Y
3/uCZCnTDPZnYhKJwu/bdzX6e7/EhaGVAGjkV3z/o2XJgmv3XtgRIbvcH+KYJnAK
mTVKRnTPj6emO0t2dSr98gGxOGVqEMxl4QavViOGN81tpUnVuFxE2vdOYuqIeLZ9
3kO5NxU7N1i5US1+HP1jA/bqDzkjJJrU0wvMTJ6BHj8SJ6VArFPO+UfxUaDqGgHk
K28z4YTh5zi1I9ht/J08NV4KYMVmz6/BeLQaFnzG/LPUqhzayUxMi9RNBb5kAfa5
rqqLacCFzaDDPzwGvEwYFFJ3t570QlJPWJ4T2tYL1+nx3tq/PnOOKeAes1JJRSsO
MzHtImoGhCWT3E80aWFDh3UBjrAl5ZqBukAt/hK0XnsgHhkw9lydrADwFGy/+dGO
CjeufmiDyx4GxilyniLB4mbt9ekyU5hkzNFG2JXR5XlYeJe1ySalVtB1iBfg6Ks4
O5Y0FkhtMuiE5MdFSOfOCzafqKhieDCmmLCjhv7X5qt6xgYC/zno9SJCwFS4lw1d
Xw+/LrKEI6pW6F8lED5En5ofRR8n9HrFAO7UDEo6WmJV158gzAQJeUrVKmr6vB1e
aj6eAfX3tBuaTV2pdkTi5IKnu3jP+KmJPiQoIjcLLK2OehE+omoVWKQc/Wnx+RVf
k+gSeHgdK8SYcydZCFX4tnAofp/GVHkr97hfC4jpiu/YDKvGOnszidK+zq7VSrsW
o+Ef9iHLCPuLZ08a1IU0hsDCFegEe2wdSxwWAVgWUpWCwOM5dlYXx6Ijr5i1PW8T
YenivPwmHAsG4BL2A3mD+SyG8bhkn4chUvtZJTk/NEqTGmOTTaJZ4gaMwwNrS0kL
SullyaAOTnlqARCbPcUFVhyTEoRuwgh9AtLs5M9JcW/6pdeuZp6U6FT1GvmomEod
adFrPVch7DI+V0f7fyueeuDyU1CBFZtceqF6m0b4sKAnEMN417mx8dNW2mAbmovv
MAij78SA4jnulreM8qlIE+gaXwOpLNM1rjfMKF0HbCj3IXPmwVrLGQPo37mm/hZN
YC5y9tKrg1O/JPB6MXmB+R+cpINF13VL1vrzyu0+zVCBj3k6wACO7w19Keql0+sQ
xnglCBEq3tpghh03a4LHIphAuLAFXtLwq9hFPFYsLL+BCwHPesInyzPoKpTSYzTN
H4Vuz+VcoDzWb+xPXSRL+H5zGYRd6Eqpe44UWprTk5cze+25GNMxC6b1yQyFXBme
xSwyKP+5yKC9vEiGPTbkl4bjgcgOUIjHbEBRxX7fDpele7XWOtizDX4X/387JUHF
7qREKdKGsTokoUV2M/wnMj39EbPktsCenfXPM5g7x5Np6PNRPlfSKC+iN+/za+Wj
eR9eIA2MR2T217dKIO/yYIQ27y1nXfhGrHEgbaVPALHz1mXS68WZvzEQPkQuC/OM
CQ78Y5REdBwhreNFo0gwEuMNa+CmqwNC988HImSkJGsYd1O4ljGwO1AhCQpAFj/X
L2HTmoFwrho1cTO8s50GUwMGZ39swQ4OESPE6T4xIUtTbpflJZrqx+bR4Vjy9dUs
kaIoQAKRLSz6Ak1k5rdTJ+xcrNDYV8/lwATg0x5TCLFcp0UaPEsuBL3LDUWCXqjG
Vkoh8lySevIGVaTvoV+uxo2lEYXARsPVg2VTgynScjjkSuz2msbPR1+XK3trkJdY
zh8pYYFvtr57KnR2ssUMYHqiV8YzJhmo94dupptVXke2dvZfeKfjmJ6SQkoPENjz
XLzmAEsWj1rEq6HUZrda8wE0L3aIMPfvMlXGY+efjnRkjTxal6zlWHD3FneNDtpp
8ZBZSc9zzpMfN7aDUENCJDNkTUjZ8LElQ17t18ld8+GADxj/s6j0wy+BtkmnY6ze
61SMxIUsNLA0N3myGUOw+U/lYNZbABs2Z3NnBmmWNdolVBuvrLXOvyvMwWr6msTj
tvHoKX8kPReuQa7mXSiLqZYY0hwRGN+tM66T8avR4sMppNZgrs1BWcaqfF/Q7yer
h9knqqfNpKSsSemGdw/9VMdW6SPIZRxs+XYoi9hew0R1qVeyZuf8DRJ4fICqw6cO
U/GKiLm/gI15xLO/SeyP+J11b1qU9O0GBjj3fI5XvVVYT9noxyTeZYWrko91cxGn
0QeEx0vmaoRft7iVtLk2WX+7A76gJfMEzfpFITNo3w7swwzNl0wrwwbjLMeujCoA
pIWzEPQkODAID9sZXCkyZd0d1G26Z6ijQOr1sz7tzFjGi6VpvyB5ASvQvAKRiwRI
wgq+9hBYT5qVJOp+0r0j6FUqGT/ussKf9RPBcnv2vQC4lB9op7u7tz2ZFBzgJSb1
UDdaP8kZG5x6Xj5+JDrSCgUBJn5mRoO+A1IIn1g00x0+7eK9jn3iazaL/LZunQLw
fWhzhQM/odN9HbC2UgXtxOhdRIsCNO4QGSS8qaoEQx/Vi2uMWce1iD7kzc8DY0jU
v5wLbeJ4CkX+2S4xjDswQsj74MPYtaOeY+O8MHpr2G5vuKKb5s8APxbgyL63tiSL
SSagwdghJAEOmnMR39LWkwGJe4y1OeiBOi0GW02FXNiuqEZBJbwoW6khXv7g3OmO
xwoIprbteICLTpjjBpnwHvefBQXiYx+3chKH8h4biSA1DzlXjy8cJKsx9yNeIPYW
5eaB8zO8eGKiwgiOoQCbYLYvZWcuSFuxjnsy5pDplqjkh1pS7GfGWb4dGfqlicET
jDdyuW2TnhxD1JQR4EsnpLzgUHiAPWSbZC8tWTVVVDPnux+H8WYgyY+hX06njAIy
PLrSuceImPDKXai7X+XefynNlcff5px7Iip8lSRoU2Ieka34+1DWrW+CCc4I9+91
3HDLaUFoxDyoNNsWZwEwCeGg5GDVQLhM7exHjHNsVoHkMFk3vov2Gy9dj1V1J9GP
KQcTfHcSpkF9zF6f/bYx9aa5noac+Iv3EiU38IGBrQE7IC6P4l4Kml1eiW+mxbnN
i0559X8OlywP6B2wMNsmQR9GP3ryRBaOhWzPF2RysQDqQJeqRts7mS0MXJ6ewE3W
x8KpSVjWxtEGPn/Qp7oCYraYAWkYcZqoykAxAKQPkW5VKxaRyxUYDfCzJcIhT10V
nYCEUjAMj4Jb1HaHueiTHw6a/Npz6jga3iBwC7c47PMNz8ZIwZLbBJq8GVMelsaL
Ycq4A/6eUhKB5hFSqui6rNPyiOAW00Va0qjBEFevJCCf56tQn9df9h+iyweup1PM
/1Vk5MUGKuausXx0hYBCGnv2H9/M/TsxE7RTI384u51kUaqCVcC3HKh//MD3YV2P
G5vRVZj0talKZOFVS1pOE0UHWR6B1ECJNDGalzXAxM0+ikZhQ36n38jJPwH8hdGB
1lrG7EQoAIFIoWLOMMHxrVyAPWccpTL7Thvog0/Etdqmjn1g52JOkxjzp/XTgIRV
9uh4Wv+1Ae5ECVQ04nXMxnHaygIUpAd9M+8ND00yDwbnlMe5hJ+abBObDk9DwRY7
bFllfc8xVN6F7ii/1kcttVtY8RIuIuzPII7FTcgrZMFLVarOydD16ecUs7DHAMla
AoCt8n0tJFkqB5LCY3CPJnlMUrtTZaWFJ/tKg7U9aDQFTIEF7yoEehyJ1QI6naSh
od/ft+F8HGGFuj0jqhjf5oJUuQOFw698k53YNa1kIEfsIM9xxMizJvjVE+JuHEJC
38ZYmSpmlaVqgAPVJN36dDIJL2JEdnV0tDHOJ5PJ5Hffb9MLgMumv5bwvTXLjBzl
2dsK9XfZQTNx5nOUrZeCkFwKnRoG7b0UJX6uh1+eGu1ePgIN4/dYDEJVi7h4lwYX
JF69iH+2p7k4oJmguHkLmppz1+1ZBpzfcmL49itN+rzcnoV4pDZD2y3ozMVCqxmz
EKmcsR+5X6Fz54Bw2KZ2gn1c7DQvbJwc2MUJbftPoDqps4ulV5J/xPLw9OkKpM0b
Q/6NV037bKWfm7NBP0KYW69VloGPCyoE6SyU1ZS+kRZjpmdmJJBBrMtN6vW1B+JN
bmT8OeqLgtVe6auFrD+EMWdbK+5NV1KKQ4pSR5r3gy4NE5MjbYXPVXeGzOzeEn6z
PAER7uukvdnw2vXY2gpyrVNZcud5iaNwLgO1949dojr+1cjcm02cRsyfatRB5M0G
mhgShH9Q4yJedpJZlE/bv+ehxuXfrJUr0owrMEawurBNzNOirN++x4XJXMkLXxcu
wzulUvWD7dCC5fLw562LK5mjZxXeo4XTVKVgUBfTvil41o7xYc1eQe+TC7sKQNh+
7yPjoa2ghgV8W5QsDVHHSyy34Po8DcJsdSzaFekM4xFS7i04e0y8ukZR9bDdKpC4
AIQnAmo6GeamK5NXEC2JlONtoL5+WlY0S+t3Os0y+hoUztdybW5h19ZqOJ4HrVQk
nJsgDmUZXgd9ktZOPqTwFIh8JEXN+P0Y+SCLOrrlXfPv8dbS4SjsS3q6HmBR7tYB
vt/2UP3MOJcViJKnfS0ea69h2RQUFws6oMNQGgQptNuRgQfjDGBFjdpbsuMdILpn
Lfs27H9Xj/RYX7ucEvk5jWIe9qRvsMQVm67JNWC28h4LhENV9jtJpDoOyjR3dcAU
UPXXw+6UNCSTeuWsXuJcYuEfxBq53vdbASPyC/Fy4SJH3dDPUv5cTXltXiNU/CVG
J59LlLNp4/keGCEyyNkYrU7Alw88shXQrGFDeOB6s4kn/AA3Pq0sJcXcc/2uBV2G
xfXLKwmXfF2aJOFfjC58VVA2JBZf6ODvwGBi2Rupckh62Zuv6mAVdQ5TF7uolItj
c+4/eCsjBBIqk0u94kj3YdGIIUwSf4BLFldnYVLSjHNGJZkh+Lv2RdDMOUbcCant
81/lnVtsFYjIGRNfbN1uHGElT0zkgGBtyj23jFoGX8+Bs4SqPHhYSyB7aBPA4dbX
rvWrK0kMYGiJKIMJIAGRreIgQWBsAUr8BIJGOG9tjQKYgZNqMbee3XwKao+Qcvp6
/sUfG6e6DEJW1Caa1g9nWant/vvBmMWIQQNp0cxEWKuPi586IG68Od8EN68JJMyN
JJg9CgWbIfEzHnnPvdSkanFRU6YK92ugTc851lrGxzFXIAJ1zgxKHONiFe3zZxEg
75TE+YU/o26yUfnJj1vWYzyzW8aGL+/MOjlpRJ5Vy+qVBmvhpL8+NHXQ++49xTf1
2T6IRvAkvXvFbAjCcxx/0iSb2nZkpM+9L5zJdsABUCmGR74Oof0zsh3kcWHiqHS4
OUHZUZ6l4iBzh4e6+2ypbTlHcEfcgVgwEdaMqNWcdQnaIYMuDKWsVnPp/FVP3N26
Calltw3V9T2qlqamIl0lKwwvEPGCU8eVMCU5sotMzMtbWNDT49PJCMhCQnASp5ab
L7bhzRT97kM0jIzKOwQ6TtqLyE8p3mDBGkuEUBeG7JOQjKLk1q1r3WTv/n0p97W/
OtWmpjMvG6jb9hkv27OSBXFplqYbrXAjbdjiSxl9RB3DdgVf5FIX0NSJkgK2XE+Y
PQW+Xl//WRw12Uzbw6g8OWUnEMMYKjBFA947BpEmX9FIMTmSDWD2tp4DUTlTUPpi
Un+RHdi3/zXDWNwWGwhBcVjRSdWSvamzOxX+C8LHnpCIHOFOfI4BMdnBe3bacC9s
dwcIK+9QkD37Dzm5c2EIFNglv13Fw+C198CLiND+/pmjmiE6DPvMGTkWJDnEWdkB
qxH91IpsVB5rMm1VlOX3TDXxCRsAslRMwNcQ60k2s3WctcoLOJx48h0e54GNaqQv
d/weIkIFFn3Hx9YAKHvOt0heiAB8VqWmcfjiXRFOuaFPKC91lD7V9aI3Psv4KO9t
l4tZV/i/6xPcgnaBE5kepHnoI6dwU9GqM2QhNHvO0WWbkArk/ukz+3X2CAMylcLR
zji4eeKeXhwQU0ssW6uoFnMbdi3Ia1j+YmHd36iGqXWY1ra69Rn3h3o2kLhKbZLg
qRJTS42SsGMy1wN7OxQOd7IwsPsuIHZE5TZHkg+Gu2q6EcPEfiS6AtpmkrRl/Woo
m2gA42+6hqe9PgIyZnKQ42NbH9LtyTe83peqMt08rk1RKwV9U+EBUC6rxq6pT8xn
by5LFX1ioKcEmxtIzmWy1mjRvUKdNQ64YCkGDm1PwmcIH3K1ZTQJsG13+MdQ6gHa
MODDILioLFGhKSOQKwrjXPCOWxMX1J1zLiPYHWME6LLUUn+3AUMLzLKQFFOyzXjv
WQlRnblLEmVaH86fTlmQ26QfHi5j5cPDCLsPdDQPLlbWKBT69sWgHuWRTVYWiuFC
O2n9r4rkAfaIB3dv6Rri8XJk5zCfAB26KHK532f22baXNhAm+QvS43eejuB24/by
JikgxhAH/jpQgglR8sZ1ZUM2I0xuwpzdHe28dG/R+ZojDxJkFM9SnFQcD/smWGJK
U3g98suGf7FmCTv5TOe4cT9ZgBjc3aAASFtc2Pi2bH3XYMSD8U7LwZWcsh76xB7Z
Zd3s3QGl6nDWQpSEk8L52GTtTIqtTplHw7CGyTY17shEOFb4FmUkJwQMm2JVxsu/
7NX+Rz1nofCf/ir+RWWPOlkGZuK4h/C8jq9YLzhmCnLlOjXCST17zI9s5hDFgwZ2
Iyl6NaEIJ5TL2cu7SPE6LY/mcKFzx7enaNdAQfVxcCcamibATq56G0M23fGTJ9Q+
5JSIME89nDcWpyJgsB0K5TBJ3n1UtljzcCNqWtjxpm8oX6rLRZbFh23PAkZZtMnv
QtAZIcZXSbLTpw1SB5W7yuhaYOKV6ya/AmzQz2UNLbEvE6Pwze0D4YR0zn3f2AD8
3XG6pK+SY+ZIcDvpz/YE1Vd9HGP4CYWyVDd1fwYOm/ZKQYIm1U5szanzLbSGvrb6
3+NPbeIgLLR3Tgf7GJ4+oXom+LMDDct4w4UZvWwFNI3zYvBhB8wZ4A4FOu2T3zgv
hLXc+BKTiNgkf1WhM9TuDqEUkg+dWn0p/CJZFNARZb6iiXxLIC+UhPBR4CYHsDnh
02kKnHY99brCg1BVuxrJqAbYCQ4UrIX5YvbaT57+tFoUT4KoxWP0w4WORSno3wbn
Icpg2SEIe9r1wztlDw6cl2cmjDLgJrmZ1ZeqEDMI3bYKEz66GsEWH4Iqk5Z+vj7X
tQ8cXg3QpQQQ0M6bbRYwc8n4Wgd6rWhws4H37l6ZU25063dEnG6VBY+K0k4QZmjC
Uh4VjIfFNcM1BBUeX2ieJfCPUbVTX2JGgVwARM/twWvUwECbNwskJYPU6I6qYzQp
dwo6LLpoDhFJAytipFecd/HLevFyoNVpi32LzYiWpktodWXpM/u7jyVhDgvzfDSh
bJeR7Fc+GAQ0zaUy8UlMnzAvhqO5hwfgSGNv1d/NuB1iJc6bIc0cEnF+trvpE8Fv
0wjky9rbUtV/Z+rh5G/vhp0MfRWN5MeYAo2Hn/JUltvmbC1PVHzxlKZo17/cJoVn
qVhvY4Sc6CNHcM/IwQyIrOcLpkWesep/mKZ9mZ1KGaoWz4UHra0Wc3RARDw7DSB/
2h8I131oLqHQZm8E3mbddaTOIzQPWmfilOWQivy7Rm4kBlKq6yq8cr45IXpanPmZ
/zi+RY/R6Hccq5vqY2SLpxpfsf34D9zgA29t+Rc41mOvX/rjaYfgAPO207nOVbG5
k5q5jD5hXNmlaApmyb7QnGRehjScw+B7cGvghidN23NN9BTEGaj/0QEw4nk1Zn3j
0FGCVTiT0d0XSFZxDTTvJPDDhxJqX+docj+2YOPmIyd/e/foN+mHSpSW/0HB3Rfr
PrZDlIbkJmMr/5b6yuoW29OwxMwDe24IxlYY3+bGNEcNBdglPiOsZLf+nE7WETD5
Lh6QzJyWfhv/pJjg3ast0+STt6NkBss61LwVNArTnpRD0daywSrhytdimPO+2ncZ
pkYyVDefnRiuLfOhLSnN6PjWZlnpUfaWQlD57WqJYfQl6ojqYhvc9NI7A9ii2nK6
TsOxe0sKpwVoF+PprV2lbx/IzRZUeBOtQbqOolZQZYwx9m01dnCTU2FqCIIkv5h8
Rn1Fn/7+dWyp/XwlYno5O48F5+nP/K7tpU01QIwP+qrJCh+c3vAJOA+oYFLTaoir
1KByiqP7njKUIczrPxMMy9pqLrPWVoxis/PV5LNe85zrKIg0JxDrO8+meKPjvkz3
bR3dkExh5fQDQpWNBgGehQox9cWpmUN/iYOU7lht3tqDX+hbsLPo+x93ZCc6bVZZ
JxDGn5dsklpYcIJru0D5e1mfQqFUdNnCAQV5WZcJB66d3LpSkiFutaFwCPeIvgAX
gg/K8dpZUfO4ibSEBbAbCQQ6zS+uL6QcLt0u2Ljp9WpCTnpjtiRrRJsuYZdJZjye
RlrAv6GlEXn0AhkNJoQuYGLD6kerqJFzR7FPBgMuAOmW9J4xVw/o0LaAK2sjJkTT
qWNTkMMDReO7YLVL1xpC7Rw0RCQv8o9YatLzqTwJT4Ob7hJ33punBLd/DPSjWOE7
aro8LkxjrisI+9fQlIshqd18PjXzbIyZditlicDkyxN2FiFgHuGWFI4Ox3ZH2Otj
HVA322+TReTAMJPfaPys2AD81kxjWJ9/lxpv3bCQX28TtAmZup6sPzw5yoXkGq/4
7af8ilXhHY6h4S8AwyYbwBcCcnTn/dHUHoGKfkvtf1c0PDpHWPQ/Essv/B47gpDe
R/bcyqLsi3ZCi7yc3cNroKBJXh1I/7CIEbWbu7+JPL7cFB7En9gcdJB2gx32Cvf2
mw9s8lajWjKuNwzMU4fpup3gAfaEYh3CKl41LMb4EzBEh3mJkNltyw24o+fNf/In
OKuIZVyub87qpzEKuPLsQbuVeZdCHE5hKYJPgkF/Cw+xgIc8KBLcu2v2pHmziOQC
11rlvaIG6lsBBmaATcwdBWt/dPuloluzw0ziVcTt4/ghyz7cO/r2ecS1Lr09PS1G
7Rgc0zUnCQyyqtS0DaQCWgvJckLVOP1YxlGVKUCjesSlYUwGzkc8Ev5Mi4y/tPNw
alDIejd0DWT9zs2n3aKZJOpXayVOUWOqOyH8W9DBoa0Re2xm4lIHodfh7w5plpVj
flpVY8Ava+wET+0aI2OU+aNGCjsL+Zihi6iOSwgL9sb9QwSa0y+G6I/JSQQ620vB
cTpBTOtAQpzbR9gvULgTmEN9mjKwMAGBi5kJRt0SPEsJBcpCJELKpoiIXoC1ILm+
udimXawUaQ7T1dPv0vvXJ+nTURHTVqBs+sdtXxbP1tBIpQqZKoQpIt4QKwhxsMdN
YmybG3P5hfrZBe/BPLhxnY7o7VkwPWBA3xfzGPDPG4ZFSQiVz6erxAQvt4MK5NYE
STXkEzS6Ne4XWKVfFiUM3Mu06f5TboYeIyv7LRC8lhLHt8bmE1i2AApCGYFCVfxV
LVFJ6y5RV0CCTjEeoHyHl9BHj7Pi4r1+OJXh/UfxQ6EVnxELBCNb98H0Cq+F0yDH
eJrzlMak7HHqGGJSzIgvd6hjEAre78rQiH5SDmacWfaIeDr9dpENW2sRj/D5ErkE
uBulrCgkfbH5K5arKZxUc6naILeHySpOouJTc5GdbF1m+Vnwel0/4bwXexya08xI
XfCk199fskB3y0uCL12Fx0T7XwaI0HCK08SGLM5OQkZ+Z6XF2xSulM1MaM2UNRFB
FT+/7Nm2WhyV3uV6zIPzr8Wkp+0B6qJNuRgfFFDDdBy/20MhBzfdMbjPF6gnu1fd
Tv1WJgOQ8h5BId4DW/mSe6ue4wYoymAz0afny9u5L+xGUyjv+veQ/1vmTfB8m8Xf
gPEuaSg95BBM/XH86cqMmDPXqr1nvmpw1+dcV8gHcIBgJoY7HucF0TmPoFZzDnCO
+Sl/4KdcWPM0Yxul3YE7ziwth4RzrQUosekWlf4Nqy/r0vRrj97aqXtx/qxfIfKo
28RzpF3tDkg+Yo3jzVK8EUCaw6fNOF05+SzQMlXjcRdcNhVjoWk9nVnKJHlePHm/
H1aw/zJASHLqJ9UIcvyPkOoDyCbsAf4PayeWbaa38wBSf2GKntcUc/1AFI+4WmlK
e/msyx7/LPe37HdMHLi3iC4vLnCPdSlNekrWzo7DzJRKzLZCe3zxTA2cTLZ3nEKU
mjKrkUTK0fZMaIquGFS6n2tDMfckI1TuX+1YfSTV2U+9QqkMZsGTm2f5Tj4k97V8
9hg0c/a5W4/kvpQvIwoHSzqNxvnYi9xKTDGd6oEftXLulXtcsRzyP0iTXQLAMoYX
Wc0m2P8jcyzGiyA28GaceMa7FGQ4WYsObQQhMZHnrDb4XVtG3Rh06btyazrW2Js4
Z5GESQ0AJ+iCHvmIYDApgSig5/IaORf1v3WR66/r+BuOWBBJ4XWxmwChn8h5NDEn
etEpb2sDsfSThK4MlxJCjL4Wkk9nub1A1lzsRMju3E9oU/I3l5ydTyhmzvSULuoy
0HbfTBERJ+eda/wjQ9E2EaDh+XlhPD0IhPT6cub812xV7g8f+2BJyZ6ZcoOZlqdQ
6Wdr3J3jzGkPzTwR2yZzu95RIyAnazlQfmWSpbFf9HoIcoIE0LJYIRGTaDkQO2NR
VNDPb1CmRjY47ztP0k5nPWqd4EBEwFLqCZY0wVh4SwZkNAuw/QncoMLEZ37iHWJl
SNReydz+XjTjje/eKOuC+Oyj2yFhCM3zz82bF0aHKaG07BDulvYK0CEKEXro1fOi
ZF9/qKX3KshpyCs5woOgsNTsNchlEWXAPCy6j9JoWpTWQhpk2eMRKcA/GDPUX2ta
7pWfswcBtpEXGUOJU6GaK0uNJ1I3WXaiWfRwGax5SiMF0lvKzde15G84/lYYkaBJ
ajUAtB6XljZEm69ds/FYGMK1bvrzM83Kkri7zItop5RS2hhKTlcmweLfKXBAb6D2
dbT8RF+rVrctCd5kJZUZw/Z7gezjuPgZfxU/1WmM2n46/7nbSn9fzZQjixSt06GW
B3219zyJm89hJdd+XAXS+2GHosM3/EIaaocU760TpK4DDciAaOwH6Ph6VAjjCulu
tf79stjqf8krJFGrmmgY2eIMhfW2fKfJF/dxBvPsErcXCR5m06R6YUE/YxbkI/gE
LwbWD+nfCEcguA5Z/UBN4iSpbejD7G1clmdgDMgGXwSRL/IKPHuvG0AsdRX7lUm5
GS9TZW9vpxxxaVqISNWdvm5J9JMGZz0q6ikBUVCF4a5R050EtfLucYOIqAdtnAUy
0la51sezQ5drS2hmvLvNdrLwpsGv+yHLiQZ0VDdZUuamGc7c0S5/UO/2mB5c9d8z
ky9/Gt5gvUD//rC2QmEkW1OXQDGbK8ZDy5mg8HaBzg6a4y6SaHxyYhSF3tlSFjAr
lGEjcFj8QdCFabnuWQPMZZ9IM3DmnEZh0wDIABU/GmbhHfK3f5E+ZOpa1v5g6ZP4
4khWIV5UzWQwYa8n9/gZEDVo+u7tswGVr2klTyH6KhcEwyrCBwzVABxyuFLZ8gMO
dg3eiYtY9OMYvqagSrNkeFMDECWv6+sY/G33KFeYeRcyjva/3RcGrN5YweGA9/rd
1L9qmjLkjo08Qxlq6+qyiwJ4ivMsKw5yNalGMXM6+TSRSlNxA52wNOeRw+mks5ST
b3SaQHCWQzwYkqWO24GYmNcJaKIIgTHwKI9r9iTBYUJU+WdhM7C5I+N2O431FabA
zUPbwDL9mmjxwb/oxpFQ+tQBX1mJGGF6I+p2iUNPPS/GSRYQ/kBWYPYaHkEMvMBk
86Wroc9aP7Qd8o1mWYjWgLdld12zJSvb33Xmd6s9r8QniioGcKg527YSyKI2kpbg
ThXIOb2ns2TG+O2hvQYextmHru5GzKlVtb2zwHmghiM6/0lqLTPCTtRVgKSGSXvS
sl/cYRx8TaR4H5OvkwAvNiP014ZHt2vjnC6XDw+O6SelYl2DPaEFkIgSmAPkPBcD
ohfx4OK8BEYHv+7AlR+hrCSNSvlk3H0h5qQoAQS73NQtRJrWydBTwN4fJ8kmQeS6
5nXTueMlC22Hghebc86dSswqPjYn3L3+y9RnZ65xAgFvM5NtQ6ECZ0QyGPMr/C7W
f+Wba8p9flKkmlC1Q9lyKvYpExF+QYWYddGV/eYp63OtUjsIwlxR2eBc/WoiBVGZ
Fs+PDa2KrKc9xC77pi00Ry+FykXNCJMUtIF/a4nJUL3jerYKPGJNrCC243Q8BXzy
xpzN5ZbPSSfUDtL9DD48b800HyG1AIKzi1y8SVj6c3Rew9yKHMBqIlkGGqEutXAI
lhIKbOrOSWLCKsLEL6eXqJkRb+JeA9AFKJHBvnZ5js/ImFisN32GwvqR7XpBczli
o7QFQPy5I8E1lhL4XoslQvpx1ybbT5KpXslC+NfowbODYW76JgKQy9Q34LW9fFbL
4BvIV5Ih8JDcUAKRVsmY94pF2nv8m+bC8OLip5X/vLjLUiuS8ukEv1xBmNxFBjXE
qa4wJVsrDpLJr4ThLTq7CmHuFWtug2c8+Ty4LgdX8cA4pm/wIaEMwj3K2I08miqu
7IWabIwmcicbVGDf7XqTeJW4YGp2i/n2ZQVYc3hCXY6kjE118z+QIIM3kw3J+o4E
r174yr2BVfIBCbGCX8UdesA93D2rscbauYNAt4ba/ehmeOpyiQoS38jSLrrb91z+
4BZh4ODMfnlASJeOsRXlDyS4AqfNxe4GkIobeh579DAXUXwAymyru3DWq+KGzawy
l64xZs3TbOLzkBoaIJljQthiZy6erZFApkSd7rm+3N+FS2CBN2bTRnc23f3ymhKk
70Vk+v74Jqca5EcMZKsbQylF42tSJqSpgV/tJntWBOSh7bW6ebtZX3Q8Fu2NOIXN
GYrcA5m34DvCiG1SIYt6+RisSjDsaPX6oXFzNtEw04idOX4wwe93vfv8hgYWDUaa
ed8hDFNMq7XzHI3bImCGXvwvKrUYUqZsaNun6HF0Ol7oSuVd16DycCM8Ay4GbkEW
Xde3NHePr0z2KpS/gVHLYNj7XcCYDl8dCRHosNDtIodFqFD8v5u6eikTa7/4NiHZ
WUlpTp3CP6mYfNfcew306QsoHGOtMz9df+OcMDHp3SWI7DTnK1qXofs645WUBFHm
wYcNNE2G9osUpuzaRryiNo2ozArJ0Ft6D+o+HD71Q6xrzycDZP+GFFTdtCBBFm01
2g/h07V5QGRNUyqwPjgaRNsfC5sNJNPG5KDei+d7I1zqIPW3lHcZwBx5ERQRxQ2h
eyfM5emQBhCluPjsNYiek72ezB2YcHWKWJW7D7boauoJ7Ma9MCzfuADkAj27ZQrY
D1eUBwHXTdhsfwZYgSa/KXsx/d12jDIXHwKQT1YcpuYfuL3I8T4uMxPSm4E8OIOU
iqSgeuSzc9l1wpKeuqmQBg8/7HzS8E8GKs2e/h9o24MTzY0ofc/UfKm9fArfyYuF
Z/T45nAOGcfUS9BvyeBSbSfPfuzNXRof//FxXjOfM4FtCh5oKc2ypmEKtC8R2x1J
cTSwu6h94jC6SX840mr6CVBDghbkohctY9y/jM1cz0z+3aJ8PUBDjKUaalDraUmR
alz7Ywwgj0LPnNJdeuFhBGnPujlUbLcHHTShT2hlaoo5EcYAz4w/L90J8HTOiPv6
/n4Rjf2dKjxdweN40uXINKXX9oHz/WNVLp323EzaZMvxaheezEByfvicXtmDhzdA
kdopxflEnB31qYm8u0lU8DCXZP0WVgx26I7RcgFTIeRNr3d31vAYY8No2EdoLAiq
9+r3X2qPar3ZodZR/smuNYa59hxBk65lOEtT/hm/AjP6RI7zg1ud1iPxWESTZgF8
U0H2gIZFo49OGq0SbhKOxhR5e0GEI5VCSExtcE6tIQ7PDNGzeENNbQgzNliGfUVI
hPaZPDi1A0LuFa2unZkvNLT9wkJ8jVcrTj8lxicNUQsFEwytgrfYlgTnRi475ggM
ytayaHCrDs/yFac684Zg9mGZoZr+tdgHzbbF3ffN/j8EqOC37l/cWIQdWWCIXlU3
U1FQsmkQrVAwm6/bxJH0G40RM6QOnchwvpSvbiZOLLrk8iLmGQ6DT+3kOlvQEvOU
eVW6s1k3MOWZ512y+3+t8+2i3cpbDZ+QJ7l9oPFFhMQWNLGKj0ux9cEnqen9sj13
6U4FfKO+jhMTi3yxvflt+7u1HVLqRzeUJNbgTSzCge2fVyTRSMCIhvHxsYdOcu3v
eAeqVQDnaM1fxRmQniJs2V27L8Cbp8V/JwtS/CnDxX1mSwYfiq/NA7MYzWO1Jj0+
E8vMucHYAcqY+MYsr9OediG3yjL5NcoweAeiGSAsGQyveNOsgLuMls7rN5+viyEO
M/geWehdvX55keS3Szki+UqviSbSrs70F8afxEBcmwZo0pK2DRVEEf5j5WGWo5rF
29jN6TaVov1RWCvZein/F7kPPJU4FaCFU4sctf6o5BCVrs8b8PB4QPQ5FaSpRFK4
R50LclMOKz2fZjiOOSdN5CjW4+PNeB9AykihC0iBcagAB+AtiG84O6GiZxpdwpqX
4afUaWWdhCaJMLSeSrhLGY04UOpS5cMYLFrXX+g/xfbykoKbRPEYoZmtRkPfL9I0
8qlecZFTk78XMkycxvbrPG8KvNN2YwzWLptgmGVI94YuslX73a94e1hSVjpsY3U4
Aemi9EEEiklX275ZhhPMWomU3LULqW0m0MrX1neg60xmciY5zs//s8Hlydt8LvtK
M7zi9x6TTKbKyuTsD09e8tk6tDFbaRYmuC6MCTSyha/wVbvGsAg9w2heUMWPUaep
NUlA+qzkAsrrBGpXshLkqU4G7nw7Oy6YC442JO5vz30N3rXhW9bp13PX/iubxJOm
0oDPfzlmhHUuCowweVj0ZuTE1ye5INkcdRpWcZxOda0YKzKKM0Bs+Um68CgYjzrk
7gOTSQWP0RJK3lCuwCDnt6Goq0/cDa19/ItlZ3b8wDGPlIEOHJosmzJfKHGPwmZL
yKj9YmVed5dYOVJBBIZRb8P8QamPvBhqV6lEH8EK7RntSyLoaq+vTflgFlhZ69hk
uWGHkXfBLm5Uq8ODMfdIV99xzDXzbF/UW1GbiZaKCmVCMY0vsmrCaN5oYnUwoVPc
C3vSs8gO/8kF/K3UFiexG9Hoabwiv7Oz6YzWw0xMCmHqAgFgjz5GTkiffA7vQU31
xJuAfSE4Pf+OdzIJsJonH+2mQBG1yI4JDLVtLuOoE/Vl71Rd4OnQHsBQu7gXyF0z
3SkeFak+bmVgbCb8c5b7r4v8wNuR/vO/fwcVRdE32WYYVlRJy50JgypmHVP92yZp
d8SfasigG+nso+5VleRXGodnNEk+OZCCZJGW4RKRQrh/nC/N0qfofTaTD4m0/eWi
6rxIc6dxhh/evPytY/EQnTjr2hNTTsCW78tUDSBfsRhjPZRsXVgT5AUfrctppm82
8rAX4TdmQBKccN2wcQWLZV14f4w5hRSNmGo0dzdcd3Mspd7CA0GCpmzTcpftfJsu
J47PXC/CGcXOISe84cIMpMaAaB1+OiJORhtbNMGMvxlt8RkPcyNrM3JA602fVb//
6JT/jYN8dq1rJW5m2MZPE2t8NnsXJ8b0xp6gRpN+eHvtWhnvtGcf+TF9z9zFxiST
PzHFjfcgoYf7A2YyWBOoIwixSb/hIhycaBR2hXDV7eUwYWKyuLxqBDLkvIxzlT/L
9JCtA3+0siWF9wyZvSRtgpXaa2G9KIyvVb68SJBNHnEQfxqdMZy0S+ZArtfMyjd7
1T7WhlQyusiQ749y4zwdMF5k04B5pBI8VWanqQQc2vm6ux7O+muzcDz/QHQZxn4o
xnyUnPZfuOWR95Q+yLtiwU+wnbl1uYoo2uYNl/f26FHMtMhBs1d4EBo7HefWcA3a
JRnm6xLgYrWyyWrvqCu3ucNzgDKRjZjB4qnlv+Muue9x62Xszr7XmZO8D+mL5dwC
fRecCwlmW9k2B690nXzxu4wA7ql/Pt9xIeyWE0zurpPodEu9cAz4cM07T8M5v8Q/
KF+K6CQ3HF7ngD3/oiYCqFoEXiUvoSvywv5bQgMMh5WrkpXGKkl7+P/JcTlj7Wd9
FenG5sTVo89LE0bEU3L2ylXmwW9cPW+XeHT9HnxBXkXrYbPRDPZyp2Qmip1dGSzj
Ve5XhQcrKuP12kgBzlHjLDFNU85Z2rY9rTo6UEEfagNmAN/hItOXe5YFFGNhlXSS
Q6OdZa41pDRdv3+9iVmAUFEMxm2Or4eOo4jC+Slr4gvIn20NWEIaenm2qg+NIgJK
dCSS/0WdW+j+asgKg+CtLfqbOnw72jLf+zQz1AFW3fh16cOpU7aH5doOznvg9Ufp
VKY97BLca8LagyX5JqXPat+409S7mbEBvVQS0Q8mzq5BkpRo57h3L26fBppIcqmf
LFe2w28V12aBTydF+179X9de2ElueYeL5jNdbEEWcgnjTZHC8KAw/Tnv/1pw3stX
NrXSXbktheNl8KAw5drwztEbQ57QoM9tFZtwR4Zs5dRQV0mSNFI8WxG6OypCg/ev
OSPKHY8Y4BfMbVV0QLUxG+G3d8MHwI1biGwJIyMDBs45qhXD+5ETgtz0nW3fxtrk
YgKmaWwsG00xklLREIpb3JP1xeteSkCoPkjmpDQw2V9/aM2qnAtsuXRIRzLqkydH
pHN3f47V2+IpPcMTmP60BXiot5/xYsWZkfLPPzwSBjgJw8V1z5NsaWgEGs+DaPvW
CIlkKQtClt02jKS7Tk48k+Ifm6vmrF0/qYlnsuHxYDDzzmXiWPxiFlQLCaqeVOE1
EqivPBc1H7MVECxTnA9PbXvkHmI9nV0wi+jg/kEuC49NwZzpdZ9VNw4jQ0FfzH8Y
9DfGoXK+cNJMBs9c90be6DBPIH7gE+i2OzWhKHdS6sP9seXHGsJGHTPAhimNxSFo
+jkOvx+TY5bjLU2qRI/Row9ntpXiQ5aMVzNh6LyKbVHg3/dmgsau5ml1b9v/aJ0u
uDVQWOGecShQ7eeKSVWHgYgs6kzvrBQbYdyo22OQy3wypFvoIDTe0yhav1y4A+8Y
IEjcZeYSjHbBiwa+JbB1dKtAxo/aS/l+DSv/g7aBW9l9hgpM75QfREGy3chVksSP
7BUBlfbl7qOcsldTSmAVmhWWBiDd3yOAT03BFEPE3RgGLqJgWyKTbUVkploKbQ7j
a80iL3CTgaOlpwb7b0jp9DsYuNwVaWOF3qDgxSI9hJYGZ7Po/QUnWI1DDD+qOvkw
gHPtxOPb36gkc4NHVdazVDPXzXg4Vkdkq2X5k+Qfy1bD2w8VvIask7yEmirFztUj
B9pPxAt7zcsy+6FCzvcA0SNY3O7xWDotHW1rJpqQEUFLypTT50x6WgwlhxAnDpY6
0pvfrO8Rv5u4bqVwFZBUH5TPJYzkq4RZY/tXpK7UCiArCS8TeUbJg5qkRd7iY6JH
JQbyHduEbNnaiJce7hhE7xbHQbtqu5eFzjvh4sxcY7SKkzzKHdsVaZVuV7SreaCU
YNW+F9PK+Jl1c5ihcLd+ZcqoekPOx9CfNHuietrVCDYev5byfdd/bi4mqOhvKzE/
K9rTX4Ps28k05oeIU4KlItvyvUrp0b08+mNatCifwQurOjo+UeFuAiH5A/JLXOqz
JMyOkcFd8IEYd3ddp3vq+jdyPFkaXwuVZUkGs1QzGiFSHsGwhnlrcqgdxq4Efc3Z
VsPEEZUxrXxnnYHmbWIZj8Yd5tNeRaj25tQNHIH+p9iickeatLAc1ObGO+46YFiD
nnCanSTx1CMF96rQ+lJJH5B45Qj6ygRUicqkrw5NE0O5qhynonhYojzMBpU2I7tL
gNMeBuQrefzJinaJncxPOGH+dpy0RBphmIRD9Czo6ILMuiAhfS1lVFaiamw8WSUK
BKsCeDCCXfLcSbAG8WfYOioNipXFQE+l4HJn5coAs+6wHJxYe1w+kxNJKD8inDQH
JUw2T7yQJ03UlSk1s3IPQL33xXVqCnZHhVq4ZwWo6lAVWUczJ5hq065jIBuA4fuY
Qf9wqOdV2FtnFUOVJ3Lu+BxalYBpA8gmaFw0WyWwi+eS9s1WlUBEzGWTzxSBeIDS
3nboL5mSRUPWE5gjNw8YOdRN2CIxMq0pF3qxowII9ox2zg8CawbNeE/m007yCjVm
k6D9GY99EwyRZbp9OE2vZtG0/+eXxXZrQd8c47D9K9JjmRpTIzCmRGiomqVZQ37K
ubkPtcHVZEqiYGosKwQ8UrLSCpUABWtoqs9OIcU4oMn+M2sI7NcfWxYxTASE3G8Q
lFszwUzdtGjAC3LjudwlGnuvRpWbt/4W+fQypkFFeNLUadH9S3JhFhepL8hcrKvM
vI60WQ4AKximXZ03nMWXUSFJ1dredpn7Cid4gAsXh1lH1o8w43wp2fEgks4Hpzri
m2McRjf0OB292AtyqLulSCMLHk6rEF3UsodzJXJIiU7nbzwAhmpA8Ej3QNFEwo5x
QpB2BpY/VJJBSC5jXOejFDsmrPk5+GfqJwtbsLbARaH4tr8bMqvMtQdGx5TjSRuy
3RDxiVMEDA9cXKwuC4kF6f1UAkA1bLfRbM2uhpO4WIiceGykqMWIft/tUX4Ww2TV
HuU8//Wlny+HwdaA0hmy/TI9J18XOs/rs8iv/xgNKftA96HrbrhjwFMAdKh0GzzS
D7cbpcuvezT03M2LJpnV+/HZQCdH6LOwB7kMiF+UNAI4kZgPkYhEjoiHn+nFUBn5
KSgDzHcSnIjYb/CovaA+UPlmO50gjrKX9IG7r53hanC1UUvyxL3BMtLgy790SbUo
H25EKwpxS5mHmlmlhN22FKq9liTJ6llDShJ8MtERMueKqW8XckrRTSdCFYXIRjg5
KJRv8UcfL5Bnq5c44OulKiBsbRepgMQaLaKQ9anciidbpkZKSxxn5wlOyGX+WPhu
kbns+u8qxaEnXBEMAiG8l3TV1Kw/8dbvNIf0cQrOPvETcrl+cQs/jwcrtzS/Wt2I
378s3rBEjC9C+EXUD7T8l8I8Yxeq5Ut8KfQtxKBneSaDlpDuykSQsfFSuklsM/1f
CKvphNF7yL7YleAA1eyPBoieXPkka7ErjH94ofCawEISyHQNYbD1LxJscXINEM/i
8nu/2SDmZhxB220nSitKK0hxSpqoJH+A/rEqpUxwJ0cs7QGAxNPsVaLXp9AfAsQx
OR5kft2jqTt525ML9eOZtlXxNR81tV4BrVEm3Dot9oyCsVEWBOfeZpTtceiZ45KM
7xcf0VVaILpZBeY35/nUvD8L6eoV8EjIJiKx0zkSihy38hiFfuPWHs3T43nTMXS5
nV20br9b7LCDl1B6c/rG9U71i1yWQ38CDG5qwPzfVz8P5HUhQMTOzNRRXqOKz3JO
+nb1rMpv/Z5c+ggkAsfxu3qOWTo/OuR8mx0hhvZb3nl07EvZSJSz7aNJEUZdIU+G
p9kXTnBmfJoxwwkgEoj7w0fRGDHktMOwDVe4KZ2jH4jVhclxZODbBQDnQJJHaN/p
yq+7ecDosGfvxbvVSERRI4VuaZRGtoWhBqmrYS4tms8lPYZCoNlkpU9mQjLwrpzK
AMHpj17BuGW6om9BTRo/Qu86ELlU0spFyOOAMRkh55HP9dz3BkfJTnZc8ZU1xM4S
9HKEc3y1piryB/3p/uSMYR380Kz5GlD6WgmVjMhnzv6W/9u5ZT77LYN81uSe9jJo
tWUXzNzgeDQfAjyH7QlNEHTBP1n/KukdbhxukouhkaxGv/407DXuC0SuvrZMXKHg
p36NQgF1kvizmFnRU0ASrN2ed/uvAICfXrCpf4zieFRbY8ZqZn33mEjFADSFr8+O
CJdo0lYTFfpqh06rXo4wzhqsfaj5I5vA7ue1ns0+z+97CPgbKoEEyLR5gdCoNA51
3Fl+KH9egF6NfizRznxUEH2KQm1/4kBxEDWH3dvgk03elmj/aDHjJYHuLLNyYM/c
UwsXEN5mph1p1vpHWkmq4iljdzZiDXjOebePnAhQf0QpnKI5P7h1dytLLQKHgJ+c
/Un6Q6uC3q64O+0zFzN7E7197YjM1xy0XBtOd5BI8PVoaRp70nVOTjp5v0gaeyYa
pzGuwzFIn5/y6drFDXX/e53/hNDB/YHo0NEd+OCQmnkz2LtE6Q7fUd+a5Z/z1K2o
zhOKj9h39Z8LdQ4kCLEE5kbt/QVsOD9ad7yRu+zPW4s6YE6yEluJ0HzzODJGnky8
3sv/EqRNDPyTsfAIpF5acdur54OatpZw4Hu1SG24mLllG7srnoBj3zPQI2fmGsgl
1rFqFioqMUqWimZn1bvnoTxIpYzjOzWDoEndMnZPOMQD19pEO8ikBqi0QuNV3mr/
wUcowrfLrxsSYGktlFItI0l57vP1Tt+Sw7smtG38uarfVIbM6s5ZSM/NFEAOk7Yg
2JgfZhlY0AhuZr9/8xuJSLco4uuwrAosuLlNn5XfJnIwLwjituj3DqMJ49gvjDTy
g9zhxWkmbg+qBNnOQjqJuE9XbA3bclKXVmgRHhi3dO4ebpND+BKiOpTwRudbU6w1
hSXuPAA7pSe7NCacywJUAoPDefEql6cxD81ygyyEc4Ii+tdgwCY+JiU/kfd8n+vc
1mEd3wPxul8cVcomemnIhyrZDUG8kP3YjhS1Q1VotauanJQssnM7SvqZoHTOnwk8
latR46+2K9RBacpxQuIUJ9gEfEYE82v4/xk9XhfUcNT/fGxVayiDuHNXCO2KnsQ8
SiUcncn45XJJz8C3m0eSiX2Xs+zKOrSmYQ+GTZ706SpoV+FJeiYHao8wQfuP+PRy
ZrMVeDWDw7PrPU8DzBtxZaylj0zPk/MYwuGIHtkgCoNuOsxAhDKB9MTUuaepD6MG
pKBSaYITMVgXHcSCAzqBsztLnHnL8ENkAlFoRDNjU3XKXCY8cTAHCdSIJP3MAs5W
NuCIcMfncS+jMq0lfNC3wCJOa2NT8C2AnyvijIro8CS8UteKbq3PoMGMf1s9A8L0
T8p4HPB1U7sTccwOe4O74PBk3wESE4vDN42P5/q1TSmh4ctSDV5oPnQJNsKmB4NO
FBQZl81JDbwfNQqoYepCG1dmKYaGPMEGEiVUl/kjSE2IP1YwGddTv56ZMCtwpcDR
m1A+us+Yn8mVC0nedpVn6K9avpIbUtZZFmz/XClU7moJTWWn5EaZHIuZhldNKue2
JtD50KgfnTRJgDKC8hCCUTDx5tDxQSFuCoKoaBkkF3Ya1jKzAKceMFj71wcbIvRO
2lI46GGpD+dntLrQ5w16xR6T8Iz7EL8L7GuFxsMXGP4q2RlP3woqM4YgqG/OCTL9
zifwYwua9vH49e89RYqp+62gV6iti5lT9DbG3viI6p/r+daOTE9irVwSF79RbZtQ
LseHQDwn7cWy2nS5tbfGYscDloNczXZ4JllG8GFp58Af0b6fI96Sj9Tud1Cf4A2o
tin98yW12lP44vhrRXsI0JfkubgA8GiRbszhK3LDTTVz00uaEDQbPmi/aXAKI3D/
Oa8dCntGbgpV2leoyQrCR7cAxypoJfLqlfWE8G0A75KIvtaY7IjPJZThdOJ7cCR/
94Ft7k/BlA++7RWLwoQdVHLAW5RVncOW1lz9zYCSr7lJIZTCXwrD0uZgSLpTgrs5
RbBAV+SuAsLurS0SAghgRdTQ+jlKU7SQJyzUb3HL6RiX0tVvIgRwiynzScbs9Og7
2PDts9c9mzxV1TLVw9SnXKdxpP0KfuKLLSR35q43CuVYsUK8S5c3JgAVLxlCDHmL
z3poDYC7j9oPz/aJk2dydz/Sud2Zbebil5XjfBF9sBF6908KdBRybH79V38tXqoH
mDiqKKrF33nx7NBkR0hv/8c0Ws/LHgLfttzy/vsN+EnlKw4a9g/HIdkUUaiCfZ+v
XoXgUFWSaFXBTMnEj7opqlVww2ZjWXWJ0zETErtvTiPpKpMgTY4RdlHM+lqePisH
88qtmHRTCBVbtlK1nIDTNierECl7ayVWK6QwyjTxsYq7FKhwBX+AJUwV6Es4FREA
i3qUqy+fzUGGAtqi53imUcHK4y/n2Kk8DkIawOd9yCJc3G6mwwImCRUOxPIs/0dA
FJwKtVryAuONivsE6RvHARYfmDNIbKbC9PqcGOuJ8FE/R8q/w8GWv71es58qrulD
wo0AxDiLjtNRshK/tqOwuBeBiCYCz1HqN9kU2KmMKQgk7aBOwcpyBIASOReBwdMp
axJnsNL23pxBzugLNzOoRxYM/pWJQ46vV6uSnstGF9o42T7oxGHfYoOEqWo0S6UR
VjigYA+YdIpilB4cDRaX3Yf8usMe3kXO/EDirMTHwz/bkI52f0HgBiNtuYHLYwum
U0m4vJTFJGZeA4Ba8YV8KrTNxZpCTjNhDD/B/sSXOV0Hembp28PYDhSgqyu7Uzkr
L1EehREpvN06q7H+6XnvQ0+zTH6gJBv5x7Sc+dftwL6vDgmnz8yVhIF3uqVoL2xj
z6ToFMtfaHjoOBzwr14jqg4Ka5JocEy5OyWUDEQuWHSuppMvnZvneyzWfsd9FTEu
FZimiRGASEnXU04vJJfeHFK3jzlNuKWm+BqBpvKDaaHgth3npdBEO9q5bk9zo/zq
H6+AHSKXqjWO2f3WwUo9Znye+AElw4TxRVcbTkND3zisQNlNwNl/rauBYRAys3r8
NaTOSPRpr8Ij+l64c1w2BGgLiYbzkx/74fWudRnzx89ZCpw3dKEasolHcfPyzmCT
eZJNXmCiUNX0oNy6eLwlzERrTJhfZlwP99XuffrX/CBJSZ5QR60tqvppUQDmPo6a
LJ2cLVHqbbPD0iIJPzjNbTZB3IhB7WBIKdsiM9k5KgwS+nSoEQxNulnNizJsqYld
jJB6G4N5y4dqN8Ngpwjq6VQ7ijkJnwqE+zZ4r+ObSOfMGe012Bf8IWoNcDK7YiK5
G2RL+j9BMl3sa9vUd4FECES+d9Ot288bNOjlVYcO7VA14g/K+pC3Wwyxm3Mnk0qo
qBL48k99diS23nZifnWWz1w/hNSYphyaMR4zjStj+5tyVp+rDXLzD2SN69/LUJk2
zXifcDjfa1VPbT2B0aRJ+7rPFw3x+H/mlrFCE7UyvZqOROPTuyMTEmej9CH0Cf00
JgH8VlDBBRgwfcrn2NWYexROYqaCose5SWaPOsp+p1E98HiPJ01CNRFdKwLlkVb1
mS0sStqhGiSidAhubGQ3QV8WhUi/7JlZqzMM9zYcJG1tAUIRCQbWxopkwP7DBwtN
ZtheQHN9qS9jg2cf47Vhs9NbjmOYclLdI4wYX1IyIPvqjWwTMUEbKBR6X6fX8cB5
wfFBwY7VbelrSKEnUCSiRSjHh3uDWzm8PqFBoUMvOVKTWNQ1uHXPrjTJe6Ufq0GG
xpsLnVKUHLwob2VjeC4aNHHWiqSwH548/X81U72m9gpzTjw9A14i14s3qcFdumRg
TuSsTqxdUIg3wsdrr9YJ8fZQsoePDLhljdeaE2x7h+DaV+hdfFff1BllARhonZbz
yVPby4JxdMDrwwJ6BpPGjpPVG6h5HNnOfzf062VazCHpAGjAxDjwD8VkVTPLzFS2
vpc2vZcd9ItwKOqMdTbRg5UK1PjFrLtJksskQ4VwvPhzTr/6PzNnLvGnM5HKVh5f
k5ttehJkDOT6dQn5pN5uvv7slSMvb4B/ZX7E/aQA5Cn96kFVw0Ii+n3UDmaHGnLf
ZdOXSOORPJNeuRLEPdsGG5hRpzjl117IZNRfzsl9B4vdxl7SnWdvEnQCDFFA/ZZ7
041Lfv2I0uluQNXlv2GALKQlPeidEbO/BNRh0gH/ZkAhamv8QE47sH+sWs0nF9Ql
Fb9Qaw34KBXSCRzaH9eMNv7Jpu3NcdKj+J6nBRLMpFvL7vOZitKB/ACK18jtLW0d
2krwGEL8nyvnY/vUnMO6sT0rp2dMzQLo9kWvVxtEsPhOZdkwuuoHRF7gCl+/Ut/w
Ws0LBivGymJeqJPX1ckziN2X832YgsbNPY+gBQ+IfbevXWZEjQ+Dbb/ppthLKPss
gARJXH/bEFEwpDBDiwahtdOxwm2GFKsawh9+T0YRI2IU5RvZLWhnUQx3XTLlh/63
tTJMFTyD1ZtwfLLewiWGSetCbYlmvrjMOHnSQasjXWcqjj6BJmCwmU7rbHkKbh96
8hXLRcR5r20ehLdjrg5hEC+cO8rGIMhaEcMo6fW+t//5HxJue1nOaGrSp5CbHXhp
Z/+Twmr0/Xi/d1NeQVXkp1S3L80+WrG1O1w+vkjCJ/xncPN0KocuDrWJap3o9h+C
nPg3sIxz7G362l0xnUkFMcHJ73aEloy0/pCskq3NvwLN+XkF9RhO9fE1S8WuAX1K
sCr4CuAfqDyzy+S2OnrVnvYlwLGh0GnvrMmlqYHCtat/mLme4r3t5SVQj23EW5kZ
t2r9VZkSdorxfgDbMcrbUyLX94P7Kk/JaVmOTOHlHMHzG3hAsOfaoRfKSR5yYe5o
ldo5rJCUCBOg36WP8PWwXnYTuEEXZIoH7tU+MvBsk9wN88AHOUoavQd5W1ZkBEcw
HTbyzAJxW07cUhtM+8hNGrBdm8Y8TNBVXHc5F4zVrwgQcrD71ve/A0/4PxFchUXa
uGbvM9z8OmBuWBgrzffKj84uQVdXLWPId0SermZN3y4HRzxXif5OOmhAPEv9Q0WX
QrAMaGZEMJ3c+g2tpHKInCF2CsfaPM/MuuMGyGUZyzw4OjLCaTKXnzyeFYjXNSIs
EuqqL8+bqQLgrFZH+fr7hRSZnQuMK00SbFKxEKg5uUHhzV1B8r+0kvZh9MJ9FWK8
wioKfWRK1z3nN65AdGteJMGfGm1EubB04tAAYtPo/pMBgO4a/g1Hg/5yscSILEJs
I0SyOZHdAKWDwjNgfQFyKmIxpo8DEgba48S/uDYpLj8/v/FR4bd/vdhCHfPG0ObJ
Qb+qgjXwv/FA08EKoUUe+/7KgJWenX+IjVyxmtJhdXPJYm5Fr9aZ+72aJej6vUb4
Xo003L7Ntoh4fVe9yrrMwzzJl0sVpKqXCU+h3T11YoMQV3/7mwrZ+jaC1AGrfji0
ugRG3BuKU5k8YqG6092vNVM34sb+ul3uXV+jflT7BmefkTMTbIg/Zhm1cwBqHtXV
hr5YgpePblcmZwYkSoWGMXFgX4K2Stomm/7XmH3hPhRHJiGUnKFDaBNPNP15NtFx
tXIyH1XAl9WqjXdsdLrjlLoBG6NejXZu9zpyXhmqyWwpTTWeGBsFttVqflpDXit6
nV8WpC/BhAztm1fM8T2MQbQXIAdQzD2hGBQkM3cIxe9CDTibagEIWst5Q5S2gYVB
xWTxSkx3+AU58eM3yzJjv/FdcQqw6pZzmHEB3I3YSvXEoFUyPmgi3hUA4Nl5aUIt
USnRWBqKaAqqn2ijxO22TFcjltp953zgv3RPDrZkQOc969xUJQ7+hv9kYlQO6xlF
9nzcI6+JCNMByHji2BuMF9Bl72jz2tcW3gpGTsAB6004PEUQTCdeeIRx8qPHg7Wq
1x+nP4+SFP5r4I82nhxgY3hnc8YBlb+WUvNrgwdxNBsCSOLvLBrSswCIAMmg1a+q
fJZuLo+tQ+WKZCxkhjZYFnlgZmZt7GAKAoSZGLU/CAxKetY9UpedrMyA/Hf1Vwi5
n+CcSqk167uU9Nn5/2URP8dDU/5dv5tFIGOnyIcSPHQsiglEEVmvjM+xGfyoiDQ8
gu6erCQAxjVofWRomWMgQW7YVAReCoCRhZInf/0Jlo6M+TSC2eykI3LmDdD2zkDg
+YgZDZP7qPhbfDal6SF8pIqo6fXJYFcNDZyxgCuuE5EyWmBKZwfr/q12eKUdhlu/
jts4b1W6gFU4snDDjLDQG78qpUYjdzYwMaN2G1PfDjc5y75Xv40kWwmY1yRiclzo
imjptFUqx/h867Z/X2xEYfIahst6OB5WadMGuPQ2WJZbRZv8v4tAm8DL98py0thh
rHLIE4GpDbLn0pKSmkJdBNypmBsnwzdgtmZa/b7yA8091v1eAiY7eN/gNlWvRA8g
oXhRg/xwGeACqGB3E+y703ihGA76gyGxuntHCxg3NcgNYO5OjcZ5HNyQPx6/SdjB
5KbTQjpxdLYbym0DBZP+2a1CZrG+ZhAdCcY/3kRMZVIPpt3ecXyK2c2P812yj+iU
hm32qsLfRyM6vzHZjcFriZatqZtPEPtAAy+3TGLZS5eI24Rsid7Huv3cs3t3vak8
jp7J8oZaArwVFHfF7Clpg6tRgNeQogszSsXwSl0Kvcwb69vcLbg/DC5RW+abSzU8
hb+6jyUA4KLZWQriuG/XHNR5xNiaoHWslWVcGFwl28Yp4OO9UyuYokp2SAreiLN8
U0AK8vAVQJ+WJvQKH1e+YWvWJG7JvMyFpO4IXy60hROx+mQ/kNcSQnVf8/X7TStn
QMbeh7r0O8P9ZrMVQS9GK28Y6pvp2XbkY37+4uhK//NSTELJofr+VxHgU2V8w1u0
YOQoyY/EH+be2MN/S+J36mpbIe9lqH8QACUGVm9YDFAC2E/84YU6D5GBxN27Su2B
AW5SdLsnI35FGleJ6649tnj6tSOOHMqGCLrD4ntV8Wk09EEMRk4Wlg19qhU4MEiS
p9+b0FbpnYM0NMQrKYKJ2aEuFNFAQOGU1ntwnuQbFJtAiDunocUUHnyaL1Kw9pxC
18nb7wdW0dCmns00nWX6rAoTnn8jYf3V1/HogY/Wi9HwnB1JWo5XOr9GIIDu/GMo
qazuP496AF4ab06FiQDXy/mmegTs0IzCaqk7FzwzG/4R1L6oxK04/JdJlQCTtxEt
wwnLhhHLis7LVyJTruKtfD0vyeLdBKkXZ7/VJgwgjdfGTFEPcki/Nv+sBCPmiLo7
UzHmTLKxJrgexi7sgs1/eXzWoDe27s08nmc5ul6x4NXBjiQHmUGx4cgW/ZHbPGCT
dtWeVnQoLdiuMW7iAQ7S3uVRklpb0UcERohgXjoP/QOI9twEzku2nO6JGI8PNvrv
k/Mjn8C58AgKm8mkC9UfKHQrEMvWdfP0b3JKOgcajoug4H1yyvK1xv27catoBv+b
JauYPctkFIhKHbuhd9w0A7NIX9g7LjZLbRqhcUnbRXumynLrd967WXBI/ELan/H3
Muqel/R3d0wDp97R9j+uJxBJjPG1VjiDfwPaeG2avKjOTEA5X8X4+4MjeetkkHZB
2fNGYM9ZDyskkcAL09SgPZ6sfn3iSh8qvpTWsBIEkGynRO3i9cqOITOP8N4jziDl
O4zv8ZI/Uh8vwETjAg1LOw04XNAYNTOl72TTLKSN3hAiA/5bMjG1UYcODZrh9BPV
njTzB4DEWlUKbzWmAPnreNpPFKibFm50N12SrD71EpniCVWnXoGrOvCO9e36NcCX
EN6/+H55Jn+lhFVsvVyy8z7YpG3JG/8KbBICIbCo9aHTTv678jkr1TbZc7Xo03Bw
e5kWuB6lyWKzBL8YisDESWqUK1EMR+FJtDNQtRiBxodCtAIplEaranIOCLdNBzel
VdrIRax/NM3zceYl+gS3fj4Tafh0NbrosQkZm2tnwuhmFgXc8AZ+RfYunFRpY3SW
34+zon10A46IICKvzv6hdMqzANQjbnhskdT4R0rCAPSbSCnBjAWypTIz/OPEw7wD
qVMb+aOSFi22DW6N3wdnDenP0RxkZvbqqAyjEYUG7K8VjBSiMyM03W39YwRXKNRQ
k8AwC7r0lVdMPN4ZvE2HohFQuCw9nXnK+SfsehDjQ2UnqKnYngbUV8x470VH5z9L
i0f+ep2vMcqGjMnfp9q44W8Q0ub2BpVqRIbYTHMJbzo7p18th/KQW6AfqxsPrhSz
hmoEG74r8YIJk7BIiHMbKrY9ZzOmCQ0zHwkPa3HeqvqCNBXcYkRCHWfS0gMxuaSO
0eGVOhX8Mao4pS3X5o0nURBCXyJaNRICx2Nw+bHdeSLFL10MwWc1r6nv5e5qd6Yv
Inc2drhZqCoUiYW4JfTaJE5qagby+T0sZXMamDr99QdyK4aXfQIysahtdgu+PF3v
9v2WTHECu4Kivt+7u3LmFD1mkp6CfNHhrHM3fgJB9MMiCAj4zOs2bXZeu/oexx1G
RSvHPM5BBxLY3aXJQ1CzPNXLeRclaTkm/yxirOwOeSdN3qY7VJzNgAohzvb0zwUK
UwngXViLd/x1cZxDfrIrZOxKYaXz/KxPSYoMo541zP6SANNFJvBD512YDZWZmrqj
lQZiBvmOqhkODM75yqTBfpSmdNdP+FuIAmfUS5O3hfRAnJ5UBtp7BZ4diNzbKTMu
1W2oEX7QPD0OyrcvGs3wIj/pyjjpU9O8Zf/HZe+hR07eJbhLUBY/wqitQDAQCFti
WzP3icn2gUvpT+BMyyw9QtNLdCNu9WOW3WPAI3BRrbGnEQM5Vw2tv7FUelLGReoZ
RPhd0o4oJSFOiD7gtBmvxjqJAm/FMFqg556ijarVq4KDU4UUsttqjQWIm2R0uQKp
YFT8OfIjPzlHuolw5HI1um3qUgQF6C0BgbXM+A+U0UexFH/84uzhB415mzf7nOC/
cCDwpuwNANrQMqqzbcNXHLYYwfjSke+B0l28q3HIW42KLG/6CyKMatxqCl1IJ0cp
2OyxG8S9uTdt6S9ebzzk6ptnNqvgQMKtTaF3nDYcAE2QJ0z8frP+vHp/dfEmOdC2
eQa3NSuxaArKgxkhjfieSHalPkb6nCt6DnSUfWUxJPvQNu3fMcvk+aZofnzMgCEq
QhXbu6TuPHokI3d8T4JBrpDCcNevfaq3xgiNr53tpgyU09WqwJltWfoEUbuxaugE
+v9Pp6LKTfMc6Avtq6c4YEkrQsqS0QFwmPUHnSjUp6ZOtG0rQFMRDuWjsgVY8r8n
dwIlvrh7lV3J3nZEMHEuTyFK3aRAMJ7DPsaW4z0ZG39DN0ILeNKCbK6tcCGYyXfr
9zGgraq5Ueo7hEjm5Ob6A3WW2Z+fEr6plEqshF1hmOFXr4fBWMuShKRJ1TjtJspD
pZI0R6KRWlxE78jJTlNVYPpbaYpvKacxUocqMwVVitV5f3hy8mwxxF90l3JF9deD
2G97pm59mEwIVuKsgeVnbU8P1+xsk4X249CogvaLCN9T+/gmCH2czF79Zg8a5qzL
2YDNwZTYg/AKSqtLzUFHShW7mTBoaX9d0Ejbz4DJnID82u08C+o1gN8azjnu1uXY
sdahzaZak3mfOONzgo9kkCOWkABjfUVziVKKEUIK8VX7omMIWkJvUcqimx8ctGbt
GEC1bqpLky5VixCNA8uZ6DmR5V2NPKxlJsp5mW9zJ532h0Pz/W70Zo6p2cR9SEuG
/E6I/uFH8/KdA34woIVjBbtRaKH/pNkmsviJpf5Um3iLf4nd75x6p3ZtjFu7tlzA
ziF5iYV2ioOw5FiqWaCHO8rAtvldVjP+VF/uivOeOTyMLd0/Xs1DHkoQYF02RsaQ
r2S6nzPe+LGFcxgGbl4vc7WbarpSkq74Yk7Q/aldD0+kmFZsHtyyco5vxMfUQIz8
TxaeLsBJmegOV+k7WiSO0A3rux8LhjtlR7txxqVUpkBBdurF/QzXT1h5iEFo80tG
+ZcZM+1Q3X4jAOyDzOsoxuKJa2buuxYHypsM/DxXCL5KaCdV14e3JJfuqxfgPUFc
8Tc0hCH5KUdEAwRmorri7oNeHIgNpl1lceDlFp/FAfMhIcKi3xUBUGbFa5oQYlVe
SZLmPFWZol+uBz3snpMA1SMoAj/JpTN+08QZkLv104Tn9EY+gfYprJ8g9kusYXWD
zLZ/wdNBqTtcE+997OlPCxM7g4kgB1lD4GlPNLquzGvasZOt+/bx1PCqnJNVa3uv
8Vp0SIz/bztlzCHiGJ9EOnQdSV8kLNaD8AraltyYHFeLKyKMcTL7se2vVouqALz1
xi0bWTnzO791o13kp+TmPWXOB7aCEj7MntmEC1zZnXRSo8+yjCZsEzoO36oHSSmn
EMB7+NJgfl6SUU9enOKOmGozVAxr0NyqGx7rBNuavRpO3kIR5T4tUJYlUi0gtnbg
8bUStLgDiuQPZmELP+2D0KLCCuGAMrI6DxyK2GvcRIIM5dQNQpqtcwxervUD0nNo
pv7WoukXTUIEooTQw8js8NUYFQ9k3TH5B0h5yfFHSa/wicZRc1VmN5QXFGOi0Q/t
UU9CUrFS6BEgnJP8sghgWGaQRGNhrQhZ2lw+TcmNl4y5jU4G7UO5z+7UCDheKgMD
rcdwzNg8rls34ZrGWz68Wszg5QYU41YaWZ1PW5wrtgqFyELJW5j7PFQmX/bg37F0
GCbH46uTltTiIaqH9iahYhXzp6nlg8NxRov9ENWfhFv3VOR7Ow5e0sI7zmHfMlnn
iXj9ZFumoAqw/vhP0lPa1Zgxr2xgQSGXMdv9a9BhRfUHpUvGk23i4/AAmbDppJ6V
5GY+pesXFAnjXIOGe5v7ViVhkdYdkJrP7NMHRLxdMe9xerBxHsZqSgEM5bG6eZK/
Cy7hQjsd2ZxyriQnYSrZNaNYVKjvKDq0Q0V7lCnJW2/97m9pyuo7EbYi7N47z2DU
FhzNH4uwi/Yzc8VFGWRwDya+7Actl3xLpTUxBdsbvhzuzk9UMm48KSLSXkvYehLZ
n43gCeCWCGjnzCf0ykfN3GPPTigoKbrr9pz+/S1uXsoMsUAI5dS283WprOTa6O6x
qB/At6YWfmyNvp6PFqBYQm7Zm7SHbiSewIXnoeg7h4Cg/mwLctNuWC4l6/Akn9ZV
/1w/Olxj41b4s6ZBpHy0IOq/6q6lnoFil2atpRz6XgoGi+4FsjtQ84Wco0QWZKhY
wk49y/vAXZjum1yy7OMQPwtItJ0vNb1uIy7lsMDVpBMwPEwGQAIgDM2t2DLOSRU9
7zSYM57GSGUPm3b1ChQbod/BzwT45zui33KagMuxbij5UwmmfXKxgu7XdIDClkaT
1lHBmJ5Tr4lC72bWYBTgpVYwiIzGjLamFSegUgxJhWxOMnWYJCMe4BHQuil+yexm
wXKNEzHQo6ZViPOLSw5gU39WTtaMYWB2E35b/m/n62EVmBsRlPpfVBReqqq4bSZK
60IghxX1XIoYYoN7PNfsB+pheypYmxZYLNdDJOutlWZwWM6UuvhrxHw009o8zwdG
sBvMFJmWiD26hUMCn+G+Qjf4/9/UOhgCeV5cfpaDivxmvZiQqbumQ10xqbReq6Oy
4KTLrVyZDBa9bQsE7jSMs7l07WnQ+o2k6is34DkoqSCP1HZ0/iy4kaU6UXUCHKaV
lNQKHJBGNnGKeL9odZqmvbhM1eO7nTaXBNQ6mTkHT1jM/X8/gx32zAX+8aBxCauO
aLLueEIG1S7CuWkN0PVkoesIg6E7QFcEZoEBD5ojR43vYsD/2P3wKt1nHW9AZA5r
5mW4a/s1/ritZ9OUv7TyjcdWwmYcDn4tFdTz63Cs+/JUnI1wGDLRXQjtvKR6ZTWA
CNA0aLqaVR20N4wcfpq7gR1K+gXb2naOozAS2q4PganVxUupfRS2Lgp5olaOIoch
5+8JLEEn/ORn9zg3jBnALEe2WB8tTAWPZwmNwgKkpuEqxuwr8Jp6q7h94KXBkB29
yjoH/P3CoTNSCpiJ/MjCqOPhRMF3ktWN7KXxBvv8JdDfNNZCYbd+Y0IVxIqvP3Rm
6CMlQyKpJOmIPdKainrI+LQguR+/YegXZ6nvr7YtKITh9Ht3qrOqMI0ZRPoXAOYf
nJnzX5jLB9LFEzOBP0GnfCCVpoyZ75fjKkcxJyQRRmSZb7cSKhXi/xtNkV9KZ6Ed
l+CbAzIO75sdfUxlZ6ogb2B7nOS5W/eiNJ7AS6+5/FqT8WEcOlpo2PPbHoROXLaF
yfFaPwsvgcljPYO/l58T6K5wB91L6vUs46NG9mUVXp9k5EiyIP+o7L+8CLRLn9Ce
ricU9cDjHB23nIFQgPtVy7UMXnZxrrMhIqUFsE7IEanHq1icdMbiUSzFulMYtjgy
esybhPagrIFRzNK4sr7u3CskXedaQt2mNNsg1As7XR1Db92eUfAfjEfADZh0NA8X
89vOb8OfPYLjSofpT5TFuBvgAsQj2FfN/WfrNsnE8zt7SQxRj76kUY5hHq4RDr+/
SMpum9ZJUbVaRTbw2Yn9QvoAqi83z9hn/m4pQgZVDw5HwxwC9wKcjNpcngM9dQAM
er+NbE3R/gWlKp/SMuadya7lYuCCVsjDIZE0c4nqlA4WHJPVgrxxvTCrwudA1POk
Xa/7oTYbNwFZHPFi8K6rEukf/jZcd2h5sdSI0h6vMH9vyV5ar/n6F0DB/WVZuiRZ
CXdt8jxWl6cIyz5j+4ow4qDBTkxt3eAXKYDlJcFzLRY0J9/EVKxEhfKeKIzhoRBi
WtOtHfz9R8GiF0Ql+1ycQO7CZ7lqRqATp26fgHHB9WCovYujHQvZPwowm9UUUIoq
3aGQdRvEl3AuY43FW+3EtlMY3xDwbuPCXKmREFroa5t1kyy4OFG7Y3qYiX27t7lA
vCUIaxzqMoCLqbBACgVlPwLnSFG5mMwtych7TJXq7N1XK8tuz3TR8XxrTYBK6uoa
J7wu02kSryD04AwYBcfb82z9InKZmK2XEhBSscBPuMVgp5MFp21O5a0XSm0s4rq7
yUIYGrlHX79TnI5hWKH0jwSUW6N1l2kW8EBnS7vGSv/1uZUgiu24QQr/7v9RVYYa
lpxAExTKP8isCzyBSeyZXF7IpBlYhzbnh0DUF5BRtF++1laEpYHhXR9v2ibSrL1B
mZSL7JghBtLqEzauoatkTYmqYkYpkObPBsxuKI76+TxwVlsu8Hev2TSDNoTmvBfO
Y1DG6vNFOoi7LaG4Al0KeFknQM3khuOFG6VxKZb3o2v//Tni2aYaBTob1/x47TVC
rlJS+bdaSBGcSd9YPzuTtpVpF94lmXTsgpv/07RcxvPhvO5HxQbctP/RrTBph8OC
vktwc7JMDXe4yqFfiTRuPhZQrlyDJ4dNFv7vbKQhfGoo+9LREyZDjx4/cxN+jWfx
LmzPWZfPbLT7jqiz9/gWi8gETQR/eIVwI0/uOKEBvU0+ELrw61sR0yJCV72SjdZ1
M5wClkEmzV57cAbC2ye09PNei4p9fF4ZV85a5Wr6Se3aschQ1j9rmgLpTuO8Mlel
KsVVzMoiQ2rnkIQWc/CXsoNHAYavUlR0bhN0h0mrcOx7Sd8CJ70x1bc8w8g1BksN
pMXF7R4kJpUbU2Sr1GqKnyWve+/ye/3Wg0bimTcczwoNWDz+gmnORFl+EoJDMmvZ
Q6wCHbyE5JuR2inhOr8ynftbeY4ODzml1GQ2ngmJ6Pvs+Y1BiIGjvpKZzkA3zeK3
doZFWHFKQ6npDYERG0kBUG9xXeG5ID99Mf82NZQJPNpdVg6gU3T9k3odntSao2AO
aB4ZhZdg+i3gxf9zxGZ2v7Xd8+q09sgf616Alxk/hSrIEiSE2IiD9lRWlYS7Alln
nrVTolYcdpK7tRIoKxvJwB7YErZt2k+435eccY+FfstwMF3G2HJsXF+8DhD2eZrd
lXmZLGqmmDiJG39nbXjQ1ZuaW+CK5k0rzAKuw8GX1ImpgAC1msIle7DMm5NEGMOM
NnbcHiiIY93be7VkY8VPFi488b8NYxDuAtaESKYCfXQ09i8O5ZkNI7A7TfiGy5X1
pAlr9SJWCtL96AgubyvwvnAwM16UVQWBcndOVMWxwRVCxwaLNkVA2XC4wQCwLOiF
qSuMQ63pXohHgK39fgDpeI3PUYnog0+pzWYMRMEm0DsaG0JhAWu/diLRC9Y2YInf
EL3TAEf5wfeze/R+JJrKSUYUjnT6tlTakMQEpO9Av5eJkR+nWLcatmgHkn+xIb9k
HyxRXZ4n14H1m2RXchWA71pmBXd5D1qNJqtR6ySlqUiNJo6epwXdm6d6nPyYJzyh
62X2FyBy3Er0PFuM7ii3PbTUP+WvXfiTU7ulH/ilnc8SSZ0wE1DNjuONkLb/0h+w
X6qZd9bvma3tCIukTsGdQxyRtzRV8F1debxt+s5dHbMtkgUB8oaelTpZuZ1Qfs0g
VtynuL7zJSFWBhA1aN+z0O2DLaIc8w6u3I7puwlck5Zpw2KOHj8LNShK7WH0l0I0
pG0ifQLwG+8V4iZ4aYgcZUreT85sTg8g2w61mF5haF7Voh2zv4NqcmQdFipjoJAi
O8i0+v0xcxMTDJxRSY6nmwJxlkNBogy8CrbqhKzHxkcNWKBAAhyLnAk2Y7+AESkx
o0tfxg4jXMWdmiD6lOHO0Z6oLs98vUaqoj1nQg/re/BNjduQO3bCRff0EsDXTLSQ
+IcFePYiPi83OeFXerjlaKdFkd7HgDY0FD+lKuFgkPbrv2QxvOzsE+Fc7UAvvPNr
3IxJ+Rofp6ZbvvpWOwAUbUL1iTirmGJMZOHQWVmDUW4zr3TLhlNV+r7Kus6nnmUi
fLdTWCZ3/fN9bXo/ZhYdnl33lFeAFQQqasg4IktnMxTkayvoCSndaCd2B+kIq/Sc
8IhcWz7lAnWH2Ji5jpt/3t6p+MzxW8xoP3WfULBwA80w+01D6dsJKpttOuvfwh5u
PNu+GWU2TjN+82R0FLmNHcH1Su3ZGpa5acjnCmnzL8HCvm9kootS0/pmgyDa+Gam
hsAxG+5k5kJCTA0eXE2ureMJ0FP1aoHpAluRvF5wJMDeUfajWKJlwlyZAfj50j0c
8A2JUlKS4qXpZd+HbuAeFPVhfz6bxGv8OmP7hJrkM3M6kiP6parQXj1mJGp6tRI/
/IAakD2rIwOz5qQ+H5lIcM3Ls8n1hzr0xRHU7s4HizqhvJviuhahoLgqPQSWHe3l
18hH+bclTB2cQ4itFqu1h4umhw+E8JbPKs7ncIjGYGM/nh0M1vlE57HuG4yQKg9Q
pnfD/Y8DeDI9R3+HbGouw8iLaDjuENIj4EJpNkiTui7linzLzV/OcFrPn2itMr1f
4uR87dCXuVi5c6TP47f7BoXyt7LSLRhu0fqspZ12WNcObm0PIMQ88/gtXzcu17ln
oC+MxkVD8DufHcCbsZMakFM6A2iDF75xH7mAaIhRdtLKR9GJAqVIpNpY9stMSrkx
/tKwPw2gyiVrK6EEqBNWdkn2RtCT0DOBI2KpfX2M0Ygcc+t3QIuLT9Hm0UCwbcfA
bd7pXr2PLFfBpnJoV1WSv7GKbz0ZhmmI7hvtL6i+/UBMAiVA7GuqS9/iIxnc4gL/
xVb1Cj46caJp8DtL8llEyzsaGLWlNqb3aKaiGLD6oNInkClahhIqN6cDlDQAki4V
WVPCm3MyLz9OjOmyNf4vU12nremPfrOr/d/rrWLlgPkJwNBQFRPhGT4gOkOBV+aW
G6LAm6GTSGN6dSfU2g4H8vUW/6gr57HHAdEQvksRhTaUsLv16SdAvJdnMtUCylSy
H9an+uvI/Rf7LLKvp+7zJBBSSA0vxWfiHlGpyjdrRKMGfg8y2lWwJ5BDDP0Cd+9S
uTCVC8Tox5lUZ0q0JhVj8dp8ykfUXztbWozTRZP6dYn8kL3zyYHLSIobcFmaHdb0
+1S10TWwePXedcJgSPXJgPfPdzEboX9cHr2SYPcGUVQQbY7hhGzX6aV4Qw2Yqo83
gEHv0QbNAQPTpLA8I4CYhKLodOJsi4FAHkwqndVxCulRH2moOD54Q3yiRnF5ZpUM
1CjnaWTfZE7aE4hRfkB0UIykywngsUPmxIE8G/LWfqZSBjrwSwxxpG/2lRHOCz88
Idm6EmOw2o8haUbjf2lqxaXf/hKNCpY6Fnh7oIocmQw5NsCVwHdVhiuvh0LpGa6k
BFnKqf/iQrElNkpTYD9WAv84bmmivofvcqQg56olSvwuB1y1UA990XlP+jww8Zaa
97WjUV+M5mf9QZI7488JJ53tmFikN7KXN5dEmwqP8DiM8vFMts1tClncjQu7T4p9
zGEz96mi+fiVH5TFZ7/vlljewYS4OufCkAN8ShVRcxo/RLXvqxYunXMS1gR5ZXWL
9nyz/WpfnQJhDPYYPkJP59y/ZCHbYwmSvTm0l39AlHLer22UIF/oaCf6iMnU1xmb
68ieX0VD42h75EzNXdZrSAln8fi8xpxFMJLsVfuEZ34WPSn5xf7plsoWvWdGEDh5
L5QGHyw/djsi5RymCaiqCNNeUFF4n+njTtvwY1v+jSaJygtpqplDSXkZV4Iucn+6
7PK4IDVBf7WH1y+JsE3NDM9RkWKp5yFBPKytoCiSVxk4pCDj1/f73nUv58YQlm0p
dWlzjEYfVUpfQjU8UCfocnmQED8ZFiJpMxFo7jqpH47DmZ/g4E1aBjCilrIjQX3T
LaLATtYijUwxBt5XWZB1lv/9faewpyVXHGLMmjOZSjhnmselzrFEwixUg+gIB2QC
JL9eXy700SigUd/OK53xkkQa77kwnN0oBz9Ycm5TmItU5Nknq/4tgvut/+4OrbYG
rfVq6tXCP8tjUTjHoJQ81BiUrqyzPU/XPtI93eMrEdzoz3Geq1sRdtlaZiBsGE1q
oDVkXO6BkXX5SA6tXRTnZBF8U2Q80q7HYwfEXR2nPIbpFpawLQojEu4leGv3vwP3
n++UbLqcN+O/gEVHA/OKKd7X7OhmQxl+mN27KwH1rUT5BZyOCD0WLCWc2Vo/Uag0
r7irS158ePqyNv6ujTyD0150zkp+6LRcMtHcRLZfyX2mt5PPV2QlLxP4lCqneGgo
J9XWLUdWox2xHDGJPklRPFVCCWN6IKp41vhCPR3tmSdvy61nU0k/FPIC/VcxYvQx
UpItTP8KoGkbH5xXzsq9X3FNyzWmeRt2pGDudHNHLKStKipGOCr3JnClpxmWlysh
4c8kQ3BBhQHG2syTECkckLwizdraStFGGghRJRSxjSiKCc7qNHoXiNkTNfcGwXwJ
5sDx3TWvDOyIXhitnO124LdsYwYDQr5SKN/3aLLJXKf6Q+xepRbz5Avf9jH0XIs8
q+r4K1On6mIpelQDzkLOCNQTqDdrYHmxRJq2cIhTd0mwENLmlXjbbe3gXnas7emV
0TFtx415DECiXZ0VjlR19KTxZCx+XLD92nq3xAp4VFTCCXuHPRJr5whv7zT0FGsZ
bMAIWgJOzQPTI4bWVu9Q42s6CiheA7nNxrzc8v2yvKV6Me/FLns/3yKcqyEdHgRo
Je6cfUTmypMpeHkfE6tfpU3+w1gvPH/lIQTMIZKsBUwOF6y4iPTAvOG9wl5o8tOg
jZCN0SMgUOIkoArM2CEXA71iYWHSVL94UpTTW3pinxF1bl2XiG7xsVez5U+UFeRo
7WMTKmJr4mKT+JmbWjTKJryPJSDayjrEr1QvBBIOPJNVviSOdBgloWr8cRguEXM1
VjJO8/KfhgNQQJUFR1G5x0xlIj5fK4phyQt+GvFc3+BgAmCrET1Q+YDZMM0RshEo
OomAzony1ziC1RtJTWgKA4eHfxusBMjjUnMdpKJGDuwx9qRMwNVOkwwrK0uZIf/c
UTrHsPacezDG1me0PSpkkQRWbMDyskceGXJyoTYwDvRl5WTgOs7dmqIz+vNMM870
KScRwQONLbGgrb2gsKyZ0bx2VNdX22bwF4oqLBsCgsqSNrPg9mAaGNRhiiSV5n/z
v/Uvuhq1NaHJcAn/2XYJsyCalacqTBxZgqar/w3a2MGLYHeZERBcRvMdRgb/qCae
g7fEeJgUok6bhHmtP2InEubZ5bOwi91+ClEnCJPM/bYTY7kUM9Ms6+RQVTjR0c5h
9hr+RQcwITUm2auLKg1Qak5xZmP2bEjyIoOO9pnc85nr0FwxvtyqudewVEG71psB
xdE2EUYdkoR+dPJXs7EAS6vGg2i7IbKNxhL/1GYxQvmDw86rU6GGMrtfCR+9Gq+o
ftvbKHEmI1ZQXUv5UfzYeBksjwRooWMhauxqQ20uc2K3jXQ40hvDELGZ/XNl7UQr
MiJenh8vwZN4oEhSS8DUULG5UgVlavuL8EoJ/ye53oVNzgRTyegJM9SO6hMUVLeO
EqOTYexseziIkoqgOblNi8ymgsmtmIbpGi9azBEV/rpya4EdSlzDZ5EqxzlqN5ou
JvBvqY4k1JPF3DqDnZC5OQX3zJKp58pQDvgkD2Zew16ivn97hHOplQt3pPug9EQV
SZW2mf4zJRMiw6GvhBkDfy0LDBWo6xhZFTfslh2FWiZNcROpU/dP0KMRJ7Swq/eE
YhCAGcHesyRD7hUadLYE9b3Vo+4/N5+QA/qHJPy5jeXnd1ocLigO/XIfxqggxMcJ
MtCnkVYBUCHs4r9jAzIhon/3NyFWZamAKD2QgLJMgSD0y8EkUtsfNlpqjPSoPzNc
4LocpjKoeJuylqRYIhNbkXAF797TwHmYRVwfjnzisMmuvJROLjEUerhRgcoRBxkp
XZQKvREp7yWk657CZ/fHVIRsJwYq6KuQTqLn2tjwZmbD74zo4uPjkB8hByq4woP/
DkiCj3nmIQz77MxsG6xZ1Aj6VsmKL4I5gbbSMuy6Wohnl5Az/zyqCQjkCtFZ5bwJ
9XKByg/HIFzp7BaxvsNA8NeLw8nq9i8I4/4Mn23SNGnT9LlDSMQaY8d89waQkTlY
Y1/nqXJglBxd+mSYr4O/Uc9RLrEpkNpwd7EwbFncMLHHVtweqny4PMm6sXzzKHIo
KY4QLg523IavodbCA5iRTaJt+jguP2niCORp0iF6/QNEV/X4eSztC43KDTT1+30Z
8JUbc3F2UVOZ8Hq8GQxz3ZGO5cbl2kTKQuez0CUA4ys20ezMYRxX0W+d6Q+fMxMV
Hbi4V5mmAFlH2qVAqsUzb85WGvUQUMu7Fpt9uf93C+JDfLkJSI2nis0N37Klb5j2
hd+vFMTRp/zKkGAqqOoZR7IDavidAh2XwVmJJ2+Kb0h3+IqJdZk7HtbIJff7ygK5
v2gW2AoBkxlqDBCWUBVQikfQJ+TpXzyV3E/iMY47eYHA7sdOI96b70legIqUwxOz
9tQkOHicz3rzlm0qAKDHZZbzyQJqvbAgrphWjWkYG4pAXsd0bdOK1H+/UibpaDhH
T6PTTI/X9Zr746jPMLH5NAfiOOPYys4FDgYGX7FcX23WAvIKUwt3l3TWZdvL6vcI
M0nCmGs3PnCCWWKMEDRC5x7+i0HZtsAlVGVnehfPAvM1sZB52cVnByXKHE9HL2N/
qrluH6SP9DWANfmDKCqH7vLhTocCXAfKF4M/PBe2Pvntyy8MD7ZL2k1I2O3Hos2x
BsJthrahLGJc2FpPuhPj3DAaD0E/B2vCaYuOjdUz3paM+FPZU2VzJ/gKh6AEbqRn
TUNm0br5JQx8zh0nLtDmc/3ScTC/RqiGYm0Upi0t7HFB+En9vciT8XvP5dgD+e5T
hJmNjWJNslZ7kvYcWOhTs+wc/ydSEWLpaC3mxdaOXYtodVFl97t9vN/szRxBubC7
Zf+vQJjsHFCsxEmGgDl9w+RrYDHk0JPM1wiNQg5Gz+oi9U8gofYVAflVg1Yy37gq
ZceYXf9FtBPbAfqwItn2Luu7jH+DXYyJVvRcTs+bvRnGg1D7rM8Faxs17IZYWhuf
H+A4NLKLETHYeMru3iYU6q+5AEl3aou/AjgvrmV8NCCaIYcaLwDZaq5Kl1/kQbfB
FZC2xfErlIeAedQiJ2rTgTqdSkYS2cZkz9u7Zf99d7aDtG76aWOEiO6jV1Tw6bBF
ABs/Ms9p3kT6ccJ3acPr3FdBfX3DM3uEaXlI7/P9F0/eJV4xVxTcmmqd/lY/bWGF
thao51TeGCEZ7iRu0X24ns/EEMKAlY9Mdao2h3kggVn4hY3eawaP9Nh7cj1cTlfI
r2X2p0ZPMRckH5wctRFFA7pJT3lM/mEQwOZNJJ+9zCK7y8fy0XJp6lLywLAViLuA
o3H1ygKVSuvu/Pw7//20EzXWAiQ7tQs23j7DbK+3/S/o5RxGVvCQaYPN6tB1SZo4
Wg7AamEhMpeoJTYwC4LcOvjAm1dOvgJLzi6fJ0HdNEsUkd1cNzN4ZftziKK1CbWZ
u1SMOC9HnZ9IkyOMW+OSs2qeKROT12NMhy/rJgFcz9Atn500fxEozrTzj6agP55I
E1UW2FBgoaCaQdhH1ZlCU2MERweYIu/xW8QL6e/HyEy6eFFrcxwUE/eleHjY7d2m
ZfyagpFPo2iye4VGHZx+g3hu2/lQGomk5dOwNi/+wdN8minsEjtvcmnBeoEy3MC/
1UApX4iCHNP8uJemBxNUKb25fDfiF88gQ6WafyPaUog6dOvq5us7TddCXHyjndJe
5on6va3Ir6t9DePITnzfbxS7OjbbgGDO1rIYx6bbB87mSIbyc7zO1lbpI8IOPM94
WOYxQd3p2AOgDVT1AIj2Q3uPGqVocMWFr9G1keWY5oisIxjaLU3xzkuXJKNpqSsZ
5irW2CAleC9agxpZOStqpxjFRETg+VOXuco63h5rpTteLEJXGcTrflz0dl6X64xZ
+ePQgmCPECyMt6/JoIUxJY7pKLSMIHR6VmT2c8NB8sbvLbm740KSAzKXttqOxgEf
M4B3lT8LuClfKSV9OIrlUaELTO4k1s/YFSZDnVBk0Xp26FwjmtOnpvv4fO2QmKlf
URXrf3QBGGagOBEBkV0DFTXOLVWldw6B4j/vt0Bt4rr3hBPvJ31k9PkW2GKcmwev
TcH0RNHU0O0h7Xy/6hjNTbQCkIfy8U58jxVvPXWX312CxFIKjPPRhujGlYt9Ku6B
hBGE3fxMh5omjy3oXMAHdpcf044XMzXOUEgFEVPzp220/vyCjipJINXiJpoV3Moe
w+/r9NiVVRF6+nJ8qnOgAeyMqUKMdE1Ouin2FfQPh3kNlBEZq4BKlHKIVap3yH4Q
3ICCLNPF5/BMycjeDZB03iMpfKXeztMCMXJGgzCQv0h2n1tA+aK/JSMOiDvWwBmT
nFdU2u6y3zcWPOsJspc4cWhBghkSnFPuQdKfns8oseVAzm0Q8W+Eb4xRDnQbmO5d
YLMP2l+oQAvWsiylp2XyWIUfUiM8IRxdFqc9NNJbBCIndWAjPpDHchvt0oynoTXX
I4CysgRKSksmr5jPOaR3JW/XrLmdzfN7UQ87QHIrwel/zRlnxQvKG/MAHOZzx9av
V6ukBgndEkRhtiLPHBMt9zNgqL/gu4KoLPDcO8fjMCdt9Dz3INV9zeT/MIUjfrm8
uSHG+kVCAfl+qExaVgCW2WFhdYR/16haFo3Q5GZMws6l5qKzGsjeZByHqKu8PLEY
+mNHfDIaPPl4EK61rHoWsV/u7Iv69IT1XRFj0j5oZxJK1mH/L1G3ZPCyRv2va8Z8
ELeVu5yraSB9n/rOCDKz3LhOIU+KnyGIcQ07kQ0V8AKWSdJwelAPbkqaWkAztbxK
b/xM7ARw5j7gILHKh7JkonHWMwrN5AeODneooj24/0iRvegu+IQF/kS1NnByQfgD
DeQJDzmIcAnCssp1DCq+mHnuEYZuMc8rPr+eD8FKLCD7x82HKH1ElTI5AwJqCyT/
ACnu1/Ck4CxwPO4titNGtGl6wDhdL9mFHXt9umyRcUOaO4dupAovZkea2m5TDTZr
lRA48sTOXKQT66+LbO+EwC+B8ozULg1RcnNYE4+p6Z65uz2xKKTw7OjusP1Yq+YR
xIrYP71o5LK+FDOzB9zOvqGgsiJIu7A8uPNtcXmfp52lUDg0/ZumFvkvareulpWw
JHhefrCEmN9uatU9sakABWiuJupu4XfKRunHobVdXwG/LVRThm56TScNjY6wjz8O
d+qvn38ox2sLqd4iazkKDM6mU3gznDiNMuHnh+ISZgQQSX/AVGYAq/anVWYqfeRt
6mXiAJWiA/4ty9VG85RKk0D2YmvK/dgkJWFxMBInvKv6rJC18xDoQxohO3nKgtT3
L1aP5qkXhdLORfFl4MDcZFE7IixlcSTnAWsmrOETZz0zcNSmkyf6JRw9z2KPYnvb
mEw+lNGDCKD5V2041tkgo/PHT+ZUkxB6uEXLGdRV/mLn59HlPuC/lgUv9dltNfcu
8lt/kznSsGQyIILkgDHpq6tzbvJyIDNUwBCx/Bhy+2flXS+/iy9X29lrUpqphN5R
F8LV0l/k06hw6rCjFMTrdP8LTaFl2D6qtSB0gY2DZIvWA/pQvSlUbppw3rzJqcoc
l7BQpWKCGWXzYPrfUTnz0XgmREgDM5xKWLCvgP3BqX1pY69G3jf8ajjjzQCLqRUA
1bpkbM/fnPk5zGr8NX4iENAnQirzGasJvvXtKoBeWYMyGt5CSczfs0bjIvQ2wcJR
pNHIP8t94z4Hs5OgSHFVwRLnBtXR5G81iMypgIqYVnrFtBsKiKt76eCgUALDald1
/iXsiZnBg7MQSCRhLgFr6iNxyu3LdvgY24EruMBEn54O+tBnQGE7Qzjjq43qBVOy
9AAbLQyoWH1Qmik59DgMZR0Icc8Hb1Y5kQNfQ59uO5J+5Avso5icXPhyhidZWFDy
j1V826PrNNoiYpw3r1/qIhy7kdpdiL9ynz8I0l6sQbmpKRDuFRl/Ef0pR5/6GmCl
jUzjI2/vC86nbFz62tNYijPkMNYa0g9pdpARg1Zqz+eN46IG+z3mWmXVo71NkaCy
Uukdsq6v8Ri1BCYmn92+v5d1TWZ/h6A0teR23oUnSDgJI5IwGyKmszNDda1sTtR1
kCaiWpY/N5viwdA9PDvWR9SNLwIPmkijdYhJzCPTQqdEVONM4U8oaAmbkcW9t8h/
g6kMDEIKO+nrKpi4UOwlXYU6RwkMLf8PPAddxnMCxIKyPkl0iCc+6IQy/lgaugBo
qjRSh+XUdJuVLcg44FLDdDucXV7VTK8lv+UFfB2a74J3KlsVaVlK0VFR5A2ZQaUc
vHKrCpbtkGNThH8SU0na4iTQz2AQVquPLa2d5qOhngr2oBvhJqJxacUQ8KNISlPy
R4iSoG34JTFDiuEXjmquingeTp0RqU97NYSIIeGK73pgaduBoetgCqoeDbEyhJCh
q3Tk+3IHNo5Ew3wP6XxKAppL/vP/EAJu3nNqxTs5Zt+5zcJ1+IXQ+GRcA7sSo+u6
SF0Wb5wbTyS65qf2gXj0AUx6zIWmEksrT4tIJVckgY5EnhvuvX2mICNMtiESzXGW
TxlLGKbdMDSY6UjURFhIQcRgxKZ8wGqZXFCIK5Y1+OmNW2leMNtTEoTqz74Cvexp
BgRilMacnTL7YCqPF+NLbGVZDki7UnzyqD+lXTLzqpQ/xpUk5U3/t7IoPmTztkoC
wH3uMmUe0ztN1M5tiwSJt+Y0+YHec5enmuf+rXtchNQz4mKMnQwVBsMH4QCsJa9w
Wx+g9IgSWfjjpPbwowbU4Vao0lntRlFX7vFaYG4tD268jDYCrCiID/Y/MOWPi1TL
t8Rws6S6KAs2aXuJ48cbeXmkrSbnacrwXv3h2eOeGuXleH8G/UgXR63XWnDI17qX
m1/PtbDxNYJ3MwiL4rzN6xNG8jZ5PDPQGp5fviepSUj2E9X0SDQiIBoTG9lCZg8w
Zuuvoi3MPpP1aOcXUfhxkqKfwf7TuVnb0Y/ftTYEuFcR21M3I6mmkip66HhRtZyU
XSChTFWRBtAlgn2tziea/I2/3cJ+HCfRNvvB5WGmuSawJTnvr5k/hKB9JLNEO6+w
mu4vmhNqnM7+NUTtmoA2JU5151IhCImP5j84w6Il6wt629GY3DanEh8C+SFJZfZ0
Uv1pwNFZjCP0wUqpYMv3dzhW6VioZTkTbCNETwURHe8j8umerAcMxPk2tmv3Qf8M
C/DjKMloIN+pcUWY0CbqtsD8gPQQpAB3ium8i//rKIFe7CCLfsT1WyYGzNHgeohc
sl3dTNlPPKo0+9E5QVrq9rFS2aZE5aah1raQj7sfj9XImf+6QO2OS0qTgR4z/uKn
bed3Gqf8Uk10d3EPO23UZK7W6ZvwmzrO6+wKHU8CkeF0GAxsh/g5WcUbOxATd2Bz
WH7bQ/naC//LU8ujB1Nnkkxtl2QGBXQCUIEchat+8aVKyo3ZwdGihB6Yl6D+T+8x
FWjlf/PZVqDSuYBYms+G49CKNaWd7KWlcbY0gS94vazIgE+PDXZRkOXfLk/4MGrK
2RaTTPOby8mPeXY6CiRGboGZbBOrQIp0mUD4h+fakiqRkA5TpAHjwSQczwZxs9nG
qDLPJlVRtGIrzgFj+1HWWTANfMI5Yb4chYZuD0JBtgwOEplf0PvwWAwqhgKD+ATZ
ykjEj6ibHuS4ol9MoL9/oOAKcmjdmK89Wp6OCkl4w4/KHnZYlQT9Knkq4gicspUN
P94Uk1sBMFGq7X8zYDPOnga0Sc7hxfa0I9R70/LsOUR1hfJrpojm6RPXEq/NM84n
GCEFIgql2DBY2XC7gIrS+KimG/LI9eULx3Uuo+HGD/NORBDhKXxmMc3Fs/IFbWso
T/of/AFWAskQ5LAPG+tOYVpOg9pdZuD50cN1BkxcnnqOL224xJ9SHgWh6nsd+Q4l
YE+0at7N717dQdvvC15QrZtKyelv3QMHpIPDLnT4L3zrQk5Fgca86gZDg98nFcYy
f+d/OHNFpVMjSj94p2wHRKSESg3xh9tAVsv3fgLeLUTHDxo+XgBOB9W1qkqYtTCq
F+w5sPt/ozIc14JNAdBRqI2rD9SIE7IcTQ2Nr7U9TF46FO/rXR4Qded4E/Ue/lGI
qsR7KqR4f4rG9VQ23qwyi2xoG5jNIFsWvK2OC+58fj5jl6cPm5qZy7vye2pizROW
7QeFsCtUHq0hDsj3PD0LVbJrNDSwRxTlbNu+rVO/rXBxkjfMvBZY7l6I+Gw+yx49
VEsIJRjW4CnH1f5+gVNn3VTrybofBkwftzzSmLv9cb8hy+D3lg/jqbLDBi7dD79P
AJhUUUhXe973BfcpwKG4rn5g0OABuztu/m5auORlyDbyq57jdW8ugPRvN0lJGpQ6
fJddbTZYcHywcO5wbMGcyWZGTL/NXM72e6B0thkfBW0FXC2qGga9tZcpMYWHGURZ
8HjZO5vFMTvTWHBsZACQEkC2urjH+6nCu+sya3dBvFEB+vlREQp5c8RU0VvBYI5s
bxsJkn7CptR9nfz21fnKfvDqSYk9Pz2e2F2ylyc+/VZY/bAern5TQd2NVFbkYszt
2ONyS0QErFN++krn5IqkQI0bcUhrU7VDVf+Eoa8yrr62XoH106FsYjaB/VzDVo/s
ZmwhjQhmxC1+OhW3f9lkaVpvz9sGle1N7zjaEGlmIIM8azatIK/eZvQrq5k+JOHA
FZpPWk2yMPAVMebVWDZgPQGWabP0+jeG+J7o9jia8mkordXjmfp0wiDhHldVr8HF
gcRQQLxi5pR6V4oDcMF7ipRe2ZpI6jq5LJPRjp3AFFWMre/cgDTHH/ZMvMJZzcrr
ZXV1YHCuX2qncifGZ4ob9Jy4B0Uz0iTpfYN+5yAe+/3rSKQpMGLQeF/DIlrvWE8Y
gYERvt64RAXij1otZOD7ijkGF7/wbRtBYRDSAOVmiah/IQhq0JxDDI1sV88dwZ8m
EPZJNmPwr0+LW6jeAt05d9QAakS7WghYNq215bTNgmEMBh7l0eE37IVCUOYOWGjp
2vip+BryHNXP1q8+xYDICy+zhaB3D4r7ulP3121/y9YuR/qnihzDUTlEe+bEk4t5
D7hjz6yuzpV9GGYW7Rkl2cT9xgAAL/ZYlhPkoamBeTGXTfENbAX9RrI1NXgNiF1b
CyPre7i0f0T1DPNFhzbfEWCiaUo9l4hONVEsg1FSTj01cmt++DgLWOgaCIypx420
K/lytJfc1ZZyfes8NOlMdNPTOPjoolZL2fMRTsh+6g2rhvt1OIy8C9wkJP3eVu0t
n1LQorhCPOxeHyv9p/fOcfKLGAZCd/P7TwdV0IBZ3lEN3xysepi/KegFfIIGZhuC
apxmOyb8mg5i+VGv4h2U11BQf16546eKr4DIxHjF3HymjVc2Z8h+xQ3V9ItDw4w2
/+7N7V33DlL2wgUM/aMzeap82yInNKpBSHqSxY/PrGKNVOG/4CwZgFmNod96IfCt
Kn5kVQXKKRRWMxTX4yfuXp1YTEs/oj2mKk8jA7VMMuGbQjEH9EjeJIY1gAmdhMim
xKYUudraviFaE9fOP93N60EEfcQMV+bRyX+IEVtxlcnImf0b182KdmdhV42JkolL
7yaitnJorC8mgp3Ab1XNMiUprKgWl3XV3uzOshlBe3DL89NyXGZi0HnMtil/3UeA
qRRESARzeNHG2L1TfBkG8CQm0/RV8sRWZe2f3AzcYRNYBmxIdswmzWOZI87qHNVW
FMx9dtc0pdRfuwAmtLzxEJKnwQcwu9RoC3Q7C/CkJMOvFoE65VU5xPPsLTeKCVDF
8vQ7muipcEB3B5Udjfh1YQbditkF/YXJOcVHvXMjzUtaUZSMmKLM+B7yDeVLsJWB
sFj4IhPKZ6YyQ8ZIS6Hji8AuoVmfVutWLlbTSy2YmmUSvQXd2R3Z7hAmLbDfq5J5
K2k8RN89lJkrYlDD2Yt/viONkKZ5nG+ErS4y1TmWPs/AjuIOL1l0LbnTom0qKJ5H
dOHnhCSg1/QeXW0LyFztO9CM+mZxxw3+lCPwcktAeraUJ/OKGm3f03lv7nTxdU3o
JNuz1nfMBSL01KR5Yt09TTwafuWWbMpZrGVKdKOA3r3XFDuv0BxGGI71i27KOPRX
1bk1KEe+kx2/K4P2YKZywXIU5Ge0mSwbNQ8NJxUzH7FJvdoqyPUhC/15+9M7rncl
1/+GHOXN8VtGqTSZHM5e8PxzX76jNrRORLTLOT3PLCsEZ5BClaf/IjHQI8mdABd5
OGemMF4DamL9vSmCLwS10U3imn2YXQjYN9Zm2M/bCiUNFOG/KiuEBRUzp4tpp5zs
XIQYpx2437qEmSAjwqE7o9Au8FXgp7+IK8p3cDp64BQWBM3dn7wpScoKbC2NG/eq
tXgXZVgyFqB1CmSJZ+fHJisiC1WPE8Bbyk/3nwFZlxpu2Kae2ZwfKAjDZLYZGJGK
/g0GxZz+tocmUdF1hyseyNSSjoutUWmMbRXGEWl/zyRlnA5IVrZymcqx9sFTM0rD
l3HyNvjEDbONJXXKFENIEnyiigG14JBeRAf3t9CI9fSYAFu/Qqoelr6fyxGlZWuM
JxH/WQpaX+POrptaWKSm6uOVrfvW6pjDvUK5epIaCJ9ZTh347vN37WyH0RWk5Wuk
VXfcZv2MytjkQnC3IOEibHocJY48IYl8TGauLy8g7A9cF/ylPHjXLPrcJPidKWTY
FqWObTsxlfkJflmGKrLbuTyWUm3EmgJIErCBSfa+PMQfyqfStao7i13rj9GH/19x
TysB9TQsQmFYWKAhkwXHBLc94rN969QeKy+2j+yL571r3fC/F7dSNLe1a/r1e5xF
Pth8109bBmfFHGdLYAMK5TVjnCR6Ir6ngb3Wj2t2V8eG5S1LqyPGA4N1+MMvbvK+
167i2orpwZWWLXeiDNvJdIGFoscN1G3zdZVbL/GH+m+5zrmWaI2zOKngS7dcr83d
MNxiW0Lauhq3LlN1g6XxjKppEVAuZGTC75TSMDW+LmbUAg5XUhwY/IsV4nq/vGkS
lbpGGma30P2DN3rj5ylVnHmu76b1xgyubeJrME/ihetkMtBV8eAuf3FYSLtR09cH
Lu6bd1idhGup5SCTjmED0xWJWu84EfqzwdCLWTGgPeDeMOA0brYOYN9aMnWEfyIS
/oz0DGNbLKvNCagh0LIrtSLL62ns1ReCMJN0tnGvR79X4ndHntzqRUl7txeoiVTS
t4SnNunGOGFuB+A/KzfAnrKQqARranoRgulULgvMOaQcmn8N4VQXMEYzgH0PBQZK
qBDRJIU0QcIK+E2Stgofwl6afCn76oAUp0P2XiRhlRRa7fbeAvPIzbAJRbD9f0zp
NgITv8RRuAn++J0w5vEPIx9s0HqmfDSeur5VpHvAwiJnNKoavN2ppgHWJAak6zDn
zT1xa/+6EYivW/OU3+9RB1TV1DL2AtCoBc/n+rA6FgScoZaJ+TJQEjzJ3maZbQQN
2K2CktzXgy6XQ6VcAlzD+DIjrrwAZngPFvkVN8oE9MiA41Oe94xIbimay4JJlQJB
dn2myW/rz2y1/KbJ1Stq+bimra32HggFSl5DwcvLThfELh8JRMvVj+FvJKInnZIC
ECKkH3Tms//ixxEyzGbroQQ4VZF28PYS6LlnAJGLspiThjFN0mq6WfiWzZ+PB6eA
4qtneag2ROrsFgjo4rJktU++yzB+O0ymAUmaN0z35p/yYuRtlzdqaZiViMVYM947
sGpd8qEqVfiXF5oPcT8tOFdoxIoFMsmnBIPsOLJfmCMqfQ08o9Rg8A0CcGaIlglf
BeY2y3BrOMGlAVxMkW2V3y1XlDlQP61hLrXvB/BJ2tPHMMW6rHeAkZIURIG5X8zX
TMlJXfB+kGy8d5WWK7cCxaj+1bREIPn/h2Jo6dx+Lp+hb0QRIC48QYEi3v0lX2kl
HGsmAMw9C2280ZgZda4ncUR+R6Ut+0usW/Mcchwln6q183m6/vsYZIFfQ4PlHYdN
4k/Hz8+tO5NJzjnEp/0Cd0FYDw21XLZ5Zg+AjS/8WuP8/asCLYsJpDb9PmgsOYY7
Fxi8kZ/wrHmc7v+bzSrO3zMajmaCBrArFdzwdD04Exz/bpn37xSIzYb6xLH8ABz2
5SZ1ghW2QUwQG/3hhj/X7mrLPGZlC3SxLPqgvE24JxElRoXjo+r4gavPstoTpVEu
Db2A+NmRrNYF3K4L2obqk60BU3LJfE3fQz6aihHR1tPneoHprvMoYWWpJuVGH3Aq
SM3y8BPjIePFWMMH+YepltJ0oSHu+1yL0Jb1Ypheia4TLI97+DLgKo+r8g7jSFWb
TGLP8XFxA8syD3XsuCcmjEGv8gnlz00VBVHlLW3LvF0b0b8Xmk5LvBViywSWSFgU
/tgGgYCZjVMhO0P7rUCWfbDjQGfO7UCcRASRO/jgVcsGm7fXPXKBzPmloJBV+W7T
HeU7q/AuRVjAJ9V8fM098b2E1z1kDaLJs9ODJSTKzXB0oIo30HSRRiP5g9Mw46Zo
ckd4NAs+POsv5MI8IUCjm5+zN6Egd7eU8+EbthXHc01eebmmAzHyr4iwlHchW1ef
rAstASiJlrjKyyWmX0kewMFYVOtS1aCz1DbWnLlOOcWQpTWrjKhlGE/AQb7SOzPh
XnfysqS+j5kL6Ak/gRTA+CDl7Cvzl08k5ANYxmkpLIH872odt3IWB4o3PVpr1IxU
eUK6qCDWlmiYOfblkwV7SLD0Bo4xPjEqJpLHj3uWGHohztxfV96Rv1N+qTAUgvmp
o1Z3bjVJ+RgB5DRkzm6aJxd3t76s1nexfS+pz58pF9+YAndsgga+muMgVwejzZfO
fr6wpJJEsBEbSU8Je92HPl2dYO48iyVwpRlzI15yKpDFtLHrtU8qEdgucT9ShHiB
sc/e4jtiBA3XiZqQ8jKe4xy6GMIT+QpJ2QJ6ruaCbMCEjMfU9E+afAiczLEN9EYz
SmYwshm9SHr4cS1VSZ7xJRXelAMoKYWsITeqkdWaoNVVWM5x5Nw/voOznp1nvHpx
fcicMTWaBCQwjp/P2q++upZ1XUVmMmeOsopHzWZNSDfmo7I9s/z1vVHALV3AEQIZ
PtDGPCrxFE0lBumI+MLgD5Tr7Cpeg4QREkKB2CorQL3KVJ+xe7DP+imKlxtEuUZo
1Puvzu4M+wUbcq7I2gxRac65J4WvO6NOayvaYZPjqz1eWrrt24gNmywVXF9owlkl
Ggny8srpGyV8hpOw5pyiUKMeHNombd3H9/SNTonaGD9GjTXlTOlIUYiHCiNBY3Hn
jwDWKXLSh1mqXaPgtHjE+8sDzqlrCJVBwQ1WrJqDH5LSOyf+qe2a72fvUI0xcZnD
iG8QAupx4Y/O5b36B36NxPLnACRK+oqs6Pz4YB73hZ82fyYc8Su8mnowz/QRBBUj
jpntIYqrrN+zpIMUx+vjciJBFBURbb6K91Ex17XzICHPX+/2dWDYnRhqfiUBmN/3
QLXgRPpf07DWHF3MID9XQan7MeBmY44QAeFVscyFGZ7JHU6d91+lWz8aF0bAob87
vKnO7XfwmWsSvD9J65Nhv3ZFfnacAM920GnxZVBKYYrx6djHOni1tDwGB0cQZuR4
BCPgCq9ywIqSaHSFTp53u5etm4OXlcFQlNuTuhJykuu8Dbuy5mB7WFMaVMnwOjGy
s+UCSLfTUAEibzGm7uj7AY1VPD0xITVS2PqapxjHi76Fd04DGUJLUcJYZA813b0R
DHwLPScAo20mtwS7HsaF8wIxZpEhq3R/nw/IwHoTz0+j9WhEYeKBK43uK6qfshOr
b+VG88e7yS8ZJWo8xkopjXw6GDxwrFvIyMLndhiMxtS3Z8+Ut8iozsdmG+8ww+ee
lN3CtgIeXKjLndTQkAj92irs0NrEh3l+vJ3VTS4MlFwRCyvTSmYJOibS3Hr7fqm6
LcEBdPUKKefbp85X2YZ6Hyeoz2xr3we02tttsfbzcTovoVDtxwnoEylc3OL0HjlB
1VQs7c67EXBSp9figHlqEjOauUF96EQmV24/StzKcNB3Yhb+gWRFblYirrBLWBiv
Tftq8QgI26JuS4AruJjM4I1dM1xdnLfpsMWOQc6/ts43RojT5T7oeorpSdFIAEtt
s89etw5oxsrFV2tRCgyCEzi/1mrgQasHclDIbGuiGvL3/fCycezT4QnDDzLWpJOo
GZsNlaw6dSeuWjlo3WIapv6LYO2Qkin2n4qId9iEkbghgDYFxrjVQeamDZmw6zrC
hlPQ5cBJcYOUgeoqcHr4qTmb+eteQJH3QsC0sM2cIBKhho9clKxHYM5itfHZRSza
LRHTuBo47RCSdgYnVRIGemBqI65MsI3/Ou2e2fDStSVZ4gpuNGiGNAckDrQTO/Z0
0rZ2PV9ApRqXKA9u9vbLXgf+ZwPQAp6WMfyMNrrYzasnRAFZOVnSRa6iKtPxzw7j
3jMdUlPgUmpPHwTeUaofgf1adhCfjoHMxXmchZB1EpPK3UusoXanMnqv0Gv3aLwG
vrF0LR1w+mzvFBlIc+I8s9pBrSiCrnfrv19wi4M1jVoC4UwohQk4QKsCkdO7I+ds
0omcE/kfNPAHuh+f1iXMIbRh2ZbrY0rfQ1qZYIHTnv6jnA+4b4jNrYNwkHM+vJfI
QPQsCuN2M4OHhHLjwz9F3pyUb3qESAkTjVeXrD4LJoqKArhs6RVSBiwMSIJhiKE7
FuwEPQUL6tqRVkPZHzCLaVdbOWaSN6GBiT9PLpUCtxeD0G/BQOpWWzdsP+cV1iCj
GSbJL0kI8NFJPcAo11XM4JzFsaMPPUt//8t5SGFFeBfw9s0DYj9GA0zZLek/NJEV
11ALPPle0jw38vvT+Toe27kL9EPnVF2cMh2cIFaewA8j5MnQgRwel/sCTsJKrdbt
x0Enu8mkP1g7fCFxBUZUTB16OBV7SRFuNxGHaA3DBdOVwFcxq/6gWq4DrRiXIii/
FShnNbjKS2VMas6DIwv1bC/wfhhhT0L2I8qQcpMAWY3BufGCqbnPqIfLPnUB0tOt
v4Xb5ZxxpOzu+UNsqd0P0HeBTHXkDwEd7qvGaIpHDzQ3lc4RdCMWxfE/w9FyBMgp
Vu3rMiFZeDq1XdpWTSpedsbPtiOc/SirkFc10vNUumRTYO/sR8aNiCdOfyJKdwLI
ezcEXabeJOBdA6/hHfHJNs06iqXRN9QK7zQjpa3l4BVB2FsSNnN7iM20vtVlGOaF
NsKE/kSZnNkje6K2+KD0PvDJCIKWocQ5zIbGr0PePg9elaaodb6E5uG8K/3mAm5g
shDKjwVSGXrV7WUHtO9JKSudQki2Dhg4oJXe1NEwDxIPSCPqEo7J7kwVVvYUeYKp
BByw40VvYMupG+aLqpbxH/gLFvpQm2mdTcRKLoHz6rTEx2NQ4iIqjsspEAUP1GnC
V9MolZ3kVRC0XaLWY19BiqcOF627pLkZHtcXYICET/NskI8pD6pRQyVly/vjtxOv
gpXD57nCAidq2A1q+eRLDhFYtXnjQx66xrv9b4Nn8AXbx/eGc79iZnY3qnLNfx84
bTgD8Jxmi1y8FQNzi+EG70UQajt2Sdp+9O1/MB/NZ+hK1h/uu7CMfbKMesiO+UVf
5IGCxb4JQQPvQj3/SnyglGFHRi2SyS4W9TsF8urdFlme1jCFPmWCBT86g5tSk3U3
q/KD0gakS7YVMdglNDrQrgxnXfPyRaJ5BFQ4PT/CSO0zpwzZ8WrZU3TzPIEj+JCy
Yp3d/rMlrBnzgbSJ2HML2bwiH+0bSfHeb9Cj+jdQwNdj9rpFjEqeQIA9z8VVK6L8
2Iqsv/t6tfurDZ6sJgVc5q84YSPLwHhRVxJ6kAHCIDO6wDzDrARRrAksk2LLl9nj
WNiJwTkWxAH0n3bw4XLLkv5vXImZQ4v13iw6y/Mov+SttQ6ImYoMCb6dhDt2eSsR
EMUYKfLtbFDi2Ctd8IKg1YASzl1KVTi6WR97jVYbKUeC5KZJQbHcIZPdaHFxwvNT
ADkBjCGtQDPMHv2No4nwSO6VHuejFvBkn8zrhLV7Q4VrndZ56XvzGDJzs0rnlxIJ
RqMzY9AGRqLueBkkIAzVnAuhwElWmJXG6blzXzZ2kebQcHFHrKnjwAEerVtZlcW/
FCDoSPwmmuqYEM86m+ywjqo+sAPmWPFLm3LUqTL6VbU2rcGVAoFsVlX9SoBM91p3
5Pd41dx4Ca6VXvY75Ck8Y7LS5d+xiGUqWgropVc2bwiFBqHch3oxor3nYuBIfFff
kpCo79ALQ5xkEyWSHCq8WMeBIr1h7ohIlIHvON0S4k9hTx/fT+3QLFshnv83FMRW
U4I8eKTqk2ZqaCq0MPGkoRQRysMnDq63ZwMks1fgxUBN5HQ1iRInSVdrBXWJbwav
m0AJEAFSDndrTdr21UjyDN1mjsaOI0JtYA9AHyYVr9M7NHHUSCgd4w4ZNGPCRcnr
Ddjy88wpqOzR37qiRdJ5S+gvi2jt5E4rOMU1dLqbYdnzPOl+PUMTBKQBSsFTtGKp
fJ2r923RBkXh1efkKSJ0thEgbRsNZPR4S9lqPTfsFX23waOpFPcziCbrhEj5wOds
jWtfRsFimLfA0mBdqCIGqZKcZwWHPnO/9C9hxazjnDwjM0H86FDblYG7lCis5xxR
6d0MwHRFMKBbtBqdbpvWLbxO4WB0Rkue0i8sbuNWCgm8JFXSAOjXIQJyieNlCfAS
h6LhhvVvUwBVQwYl7rtDodsrhRVOSyQh6wHIJalu5MKUX4NOtKzpOmKleuTBhKp1
CGeEE43F260KAVvpDXLQV6W2KOwzn0TuUvig/YUuIMfweDlWyYrTj9vp8BGD+Vmq
BCQ6+Tam8tC3vqaAe+NpzOnwJ2MHK7fu6d+OXWsDGBgP20mWG8tlRyzy8A7p5RvX
iYx/n4t0+i7wlly52tjHHvDueRzLbp6Fw4k8EfFgob0lB7OIlJ4xb+qWqpSi3GZU
0e8n1k+tRCDDFSt26w9+IxDt44zebTNeWjcaDRDL2Xgty/M+AP3dZbCJb6QsTY/f
nxyxNq4ivfEph7C4nLaDoW5aUng6mgiev5/sx5E7tMumkQQpWJLotGRaChJPdqRP
d3M9zf5zWK4GR53IHB+k13mKUNV4fDiGv8F97T77YyLdupZE14slZp5nk4gkpG63
u/5EZ1bjbLgwBqUq8pZ33T49xmaouQM4SBf6TYCP6zp/KgFxjug6z/tG4eE1EtMe
VlrizNCgZ88o/cWe+BnPCCNg6oyID3f/aU9Y9W9RFOh078IU5TjwIOEIMNXBs6b0
Z2l7Xz9YGBVNk6cGW7fDGCZkAz0CmTB3FTFrIArUHLOO7hrHgmtjIzFurMDLEdst
SX0DMAN4PBMw1JYiiswshMYe0iduvU9Xe8slHwy3Vrb1gb6Qkhc994rMchJA2OC3
HoCvVqbRkl/nNPgkHZghJ+xBhDThfAS+Nimk7M4PxxPiM2G45kwm52teX9XB1MHK
jnfWUTPcsMFUlYDwVFCBOoRpjnv9g+5k4Aix3hV7rj9ysV0azeUes9AjfQCQjSTJ
c7GBXcX01vkJAAdoz9WQh9K28Ud7mYtjV9AqAs/+V2YN/eK5Qo6pmkbG68YlnOrw
M/3DLHQvXYoIOuxSRH0Visv1boGZ3+xi58PpPYBg/DZPSm1+CHd9+8R1QPiRo2G4
OP+nHlaOl4j4SgUoAB9ThoxJrUHeNOxXkjs34FJE2NjPui9hXpdfxALLulh+5TlM
KGdrI0368ZBt4J5s9Gf6gwG0Tj+3EVk71A4N3cYDmZ+bk3QdOpXjSOuA9n/msSNs
WFSofAs4B5QwGA0dljbqnmjtH3MzbH5Y7SebBHutZIv8CY5LTup2k/Gquw+rLsTB
u9YzS3PjBQgMRumtvfeQMzOfQ5NW38P0e0ng7Q8sByoPEJdwVr9Rd58kgJyp7Ibp
1j0Rdzy430E777rllrdGovFMwDOh/1KjxK6J92k1JQ+6FLr4ZKCwv+XYy1RomZv7
mICBrjhTRQftldp37KRhBgGNH2il3jKgH5shA5euuIfU6Y31sTIk+VpwlWls5dOj
VsmPIGImuuHf2iwPlm7PgXHqtydedeQNFkrDn4xkkBTouOmSny5E4HlRpwJiyxtL
clIhtZRcHWVa2fYm4eshUU07/kvkD/+IryTk2zT2JsdpdewLaej0+lWQAdrjiBPV
GYcEUVW7qLG0hzSFYUthwvkJlrtoy9Fp6nCOUvkIiaxlJnJa4gKtaUAaTUi/zvQN
ie8s/9qGGUEjtd63lMIGxz06xxr/FerwHgzbnMekenmbVE1RlZdi/hO4jQY93Vgp
QUsHssVlGAXiWwL7fwhbfwWXz0TOQJqEEDLA6rT6jLOB062kuqYF18B4I1iEIENN
DdmVs/21/p938JprYIj/iruq/qC8qjfrC0Bay5MZ3pMwlYz1E0OouAxQG0McMViR
MEHcMJUYg+0SuBx1TdEFbweHlqsXOJHL0SKSuFq0Oqly2zYaovUffYNBqFxtJNw8
ABDbmLmmeJDCCYrlqxpLtO/Nxu8Gcp8SRH8/HtL/OtGLOe1GabHWXo0FNLsimXNY
KDV2FSdzSxAvG7Wvkkuf1gz/cDi3FpRZ6sQgDskF0cJLnwG5sE57usTw+HeHMXAe
NSnw9ciVhJh+UvMZgYdNWW33SkbnAR3CDpnjTXLnJj3FR257bHM/QGgENewJG2Py
uRPx8TP2h8h6570YiYswLA7ronGwJyU8aj8E2Rtb4yYWk6uJSHOUhGV+VKQhOa3L
1PO/WgkWt2pXpHb4D4g+xwYNhgL2J90er24sMrnnvCGKUw01Y0fi2bmM3v0vZuUU
WNfxmm7hPxT1s1U4RE0+WDSbQAsz+KSBIs+GrcuTq0rjZp7GTWU11x8CDbVp/mkh
cdGxUxEYr6MIaOqNo3roI90FlTSDZMT0t88/2/cC2RSJBolsTccuWnx+JDvHFDvK
PxMXYDGify9ZrLqHCQfSAW+aUv2Md4L1REvZCmS2xKPe8v9Jto4vVG7qAu0AUeQp
Y3Xi40xc83ADlQpJiOS8zwrhdLHyDQb5s2M/ArwGV/5FybPkzgEhE5Rv2rtNfybW
0k6v0Vz719Dig8spY4XmrHmLv0Q3sEW5zVJxDM2LLSbJS5xto3L5tsJ4I+hu/9/x
NZQ5I6JAVJetOUdlJBWWKh1mCNyVQh/ogYWUXiPX+yoarhXWlgj3OsBd4Cxa/zd1
EOvCWdN72z7AI8hlH+3BSJ9c2SJ0O69TsQ91Y1CO+dHguIm4iaUUXS5/nHwlx4Sl
detReE4fbHqxcctLDI62UcuRP1WSzFwkhgDGcyjtKhxs8rdrlSrKlVN1GS7wARc6
XJD/p2h6I4EDLX0RWyIFt9UakxeiZXGJHAJQKqXYLRC5ghvH2UwVYLdU1pQ4PdhH
9KwOdP1sXkmBU89k/LekjS/+mvgrVLFQheVBIXXareZta91fgNfAUo1HoyI2jejP
cqILF6vmdrKQN1Ikbl/WzEgeSfgoWkeNEqXv4P8yL//SB09qOZI1v31wWYl6yPR7
q2UDMhxYWqZJNMLGfIuPcDbZ8FPpv/ZOJE29zZzMIu98zyNeY8Kwy7OJoSBxtsIv
gKtmN5vxfxnvb9bYzm1PWhBAybAKg0EzA8o/Ldfh+s5PM3IuauHfp9zU2MK9HW0D
bP/cZqgL13+LhK+ZWn83ljfUOn9FTMcm4wfbrQ1SSIGhjZs2EHNVoXqIHLHAg48R
KBhBVPtsFV76ilHDQg2mhD70jqLEJ1Td8kLz0mf3NJGK4OAKk180ocooBunIHnM8
NLh70sAGJoZRtukSi55n9XZsOb5wiYccHIEFVYdGHI7Af+eLZU1VodffbA0bmreJ
Osjb5psiCOCDLCGmAhS5k5IAL6WSUur9KQOWnlf2UBhIS9wQ1VrFZ0OjQVWX3jfg
OORv7lsHrwa0RwS5KtUPwBYrkbTwRMtbfg/k1MZ8fkuOlk9LutvYYHo5zYzjN7kx
OsdgSnvi5j7XFu7qi+oSqER7uL7rhpdLU1Y83vjbq1whBIBgUgbVCLxGn/JTCe2b
KcyboTgGil14ZZcOHdl9BByAIzd+D0nkNlIjX3Ad3DF2WlUuBxCuBK1yTPJUxsiJ
zaiP2lbt+xczi1XBkAbMVghHzjGdbJ+SPr9rXZVhTVr6Yi/j33mBGyr/fKKZVc4s
eGpo9cm2tAy3MUuDaX2a5ovSEDFrXy4TGC7Q+rzrQLLOR2KrhR2LScbfwSe3vL8R
+YK9byfipML81HX4ywCaqcat5WyR8tbcb6nrQVRKnhHW8jn7CIw9e92pbUDHng+Z
lxHgQizryCT59uRHmbR09oAiUaiexjDN5K1yGq2PEQGSHwLCboWRrbj1GXGdl4ss
8MSDNB6r8vi3G7SGAQROArnhFsnB3rRzbPPhAAEbMTUjJRhyhpBGURedwPBE2M4c
j49MrlZgbtHLtbdLNZssdkGLiNyftvrS6gharsr52HYz9yWkKEvwBAZeKrUZYVAI
2zlMAljhf27su/I3u1TUWPueaDY2h2Xksyr/o6c4d0wI3gGEGBe5jOqFveN0AmkS
GSfJrnO/q4NdXVDbmxMZzw1CXxZhyAR6Tq1semOGr/S0dS59wWhorzN+0y8R9y7I
Xh8L9AxKFwHqtDpG0GcMeutAcRfikEuja4VPK7dm7O4O2jNAExuv3jAAbfGGtN4s
nGBwzMSSir46bP5pSu6YtyURo2alGA+PRGN+uJmQT7+hv942S7DZLXSHbqi5/3a8
9T6oPv5Q1lnC+Pn//yHJrwzBShLPpoGTscEnMl9MJQ/0+4h3obLj8ekPvvdHRMjl
LxlMkrV7UMkj2GPC+etPhOMv6jL2A84RbjKqPfc8HeQDR8xaXsyOZ7BUTY4zZhp0
/R2WGGfg5JPIYxQZnx1oFWEuI+1FFFKL0e9XDymHKU8V6WFRUI6bPVO3DFt7pN9D
Bi0mIJ5Nqm2lQF3TZe+cKmz5tWdJccbeTVjN9Q5IoBuBLnjc51fBeyFioKrp9MWa
f/I9QLdaoI77Jy/CyKiTOktK6jJl8ITdFeU+Dld/3gjFR7MgGx/1cGsE/yzkDlZ5
1Sgdcf/Gg2GzGoEcMqG97kzVq8BdxIunIts76I+PJBFQAtkynLAYjxmDacrsVW55
PhWAD87I7loentW10DL8uYipwzS9iib5HJldqzeSTwrrR8O1TU4KUrFBG11URO2l
2WhqBd23TTXNtv5FTHt0CN8gqbtvnYyrxxbk6wltvQ5s+xeuB9s6I4ld16CsqeDd
zzgJ3UNxLgGccPEDuWSqSC24BOhTkT0FcBENySRoqoxUneqA+FQbVVFeH4U2Hbo7
9KUV/jjmMHhEtI5biqYWoLYQxA5FDDOus9II+XeZURxJ0Vx5RZ9+Mu9R94ceSjky
zN4WN5tzZ7eBquWsT6axBhmElBSf4md8knHBEwtMFq+LGtL7e9+JlG6uJaQO7mXr
DR9OmmvldDQqmYOik2uDWpbVhVJ7/NcLU2lJIkEC4xRxfHBLTmfLl86KAT9BR0Nv
XVWVq32X6tieSXhJNeGCxdkZ9HFCqJaMg8o3rmhoC0ZI4gRW8kUIwj3GrGbpo1QG
JJfjE/pUdusn/4k27zSAb0X8fO0+eAsXa0sHiTZEmYgPJmJipDdCsUSC5Uzp23SZ
37QyqZrEgDD/ECLnf0cLfQ2PsHXvvlROVHKWsFMJSYN8T5wuflBH5PSR1YfPQQ5o
9V2WlJ9uyxGqsw/GHHlE4+nGWUzd2FH1LMuQ2ScSDabRc07OgAImsLAZpe/s9xpn
77B8gZZ4wlHnz2dehM81P92I66+j+ckLADSa2YNogorW207J1N5S8uObTBOnES+f
NozEdN260zGc65JuSaqDWCXAZZ4FPVK6uWkNAo84wsNd3lLwhA2G0d4244tass0D
qCIlXFLPFWHksWxfbHaxaM6sfHYsJgW0zUqsLHUjMK4cciQihqyflBjHyCbx4HQs
eAhPW+I++TnZLsQYBYigaPfSy1DfSDihTmwGyc4mRVdpQdjW+v6qJxVVvSvjt8i5
Cw9RkfHImWPhjpu+0bertgsZzPjP45bPJ0RVDmCAvKus1coff3H10llGI/EgfWfQ
622iBEcSyCu5fgWStWfMmy4pdMNc+ol4oR1hXxN+tSApQs9Ocoqf+e4NBGtJYSlw
LBZi2cFt/+SuoB3oKFMqLSHM++rYkbwWMg5/E421t9hCzbuBV0UQIWwbcHpFCKzt
oNRBAER6jjPeJh0yIGLbp5mKCVE2Tbw/yds4I8Kn+PIOqeHHXsTwE+fHKBpPKk7I
BcED5wruQFUfgScwMurFCH/D624JXGChR3u3LqeBq1c6/gj/ktCxtawVWwhHig6A
Ir8jhquDlwm4RD+HA2AXehv6RonNGVhhrnOXiyDGYFC0LDYecz4hoPHcyQ7u57Cw
xOnVFl8Ca5g61+G+XnqymWt8IN+gDabqLbtnnKyxx0GP3N1nccNQHlWCqOSqnIqW
eomjdKLB/OneRGtd4Qu+eqT0esXv0KBcxgkuSa5goF/e0FJqblzusQjWBtjxoa53
FnKemFwmK44Bhy3pExPSL2cjtFfQ3ZmkKUrbUalWsWMZIX7wB6tOvpLFy4lHsT1N
7WESB6q8MddsdlwUjQ7XqjlEPncD+v33ErYbRon7xQAvDNKWxDR/Cw1BZeCqvPxh
8wQvi4RxOxESMVMrBnJIaVXU0HuTK/Gs04OWo9e21ExuiQ3zHLYWAZcfMU4uauta
1cLxEB2/M5lmI76YdtIdpRghu/+HPlsvFhs6SeZG1ac3tf3ECkI02o2WYcb4vwHR
1Xcfs7lpbQubKqFTDp6nT1pCESiUN2y6v1A4kSwsYAPHbFKUMe5WIo9pG613t0SO
Bb3xVku5bUhumLs5jo9n8qvc7HbVeB6d1hTkQ5bg7XvDSwyRG4bU3HDBqGP0cONe
VT/5uiG4gaDyYHZKcgpW5rxIDdnR6XGQO4UK3YxLhCbNnZlRvmJise1eJqmmgtJD
E522roNhzuHUDpH+kF34KqH4G4IcW+t51GevcofreXDCUGK9Olz6RDLUlzkTE+jP
kmD854E8ozcghlcNZkNClAdKqOFiwHLrM4aNiSqc1WCmy+6LnGQV6M99LLNKtVJP
niIECim3WvNj0oS4xnjKLgQUuODJky0jOP81VInMRrs2tqHR3MqG5/A6RucmK+Bm
ba+GkPBiBpODykDe97pwPwPzicnPgnFjmB9wuB8q0zpcfDxtSnU0TDqLsFlpDVi9
nyD3TqrY2MvVRgb9N/q+Oq4rFzTKe37Ycsg/z3m1x7I/U/x0ZggGcpNCRxF/hn3G
Q8RXKD8UpV8nA55IsDYq+ghtgKzt9P9crxLJpboP7tPB2QVWWMlfZ/7ouoKYxTrk
kghOWRcxiLNPARuXaUgxb83jg36ZM17D12wACq4a2tZ/iiXR/ab0bkU1P5w8hidp
638dUtwSxSh7k1CxpEd1P77A9zHYDKSTGH5akZY1wJhetXq7s5EAOljeJ08F5Roy
r023/U4qB9LcQN6G527OrRGLRebyt7f4KG6RwuNDqdigQU/cu8V2jvRjKmmduX0V
qo+e0qwi/yiv25jYoYr5gq3z3y6gzD8HJalRFEz12zMM1Mt96z61Bzrv5w6T4ejj
1kIMl548VlY6uFESxRcLyVW+VNYmA4tgRTtv/fzjaEsHgfNhS5nQ9jSR+j1bNW36
Wv+uc83k6u8FbuXWzGl3xctJ9+wvq6QK2373yrydWi1e8Niwd2xZxt3pZyJDcRwA
UpfMEo52v6lxbiqSRuEtIeDMnwTE++H18lW+1BsuvgIYda632QQbNpTF4uYqF1PA
hDaqULelFDmGyjZ4Htv2fHXOeJJhI/hzLPnvWMkzr519hli1h8N3AKQVT+k1upPi
jRtDtnmlAZ6lKJ6JVKHz28FfpC0axsidB0uz+ISami79GN9b5f8M+rn65DIWWpxv
wOYrj4c6zYH3+G0sTK78eqgPL5TRMThwOUd1s9Y7EIe8wlevEo++3O/Qaegs9kox
Sfwu1OFwbnh37LQGYq329LATV31ye/U8tUOm6h7yDAuZYItTZrxb0gAU9u1zKw38
2sYxv7Z0N886HFyiJFQ7jPCzyPF5YSqPAUBRbwbVjlThjHiU9uKlsvZpLMuBXfV3
xYXxrpcfCl85UiRh1w2m7n3/zi+s7bIo9whHMd7WY3cdHK5xxeJd6DI8m1WmOtSU
pqIuHAGqBdUyVdlVkJyc9I8Y4AIY6XrbFAkuKkN2l9yMMipGx3XA4TAkYg6wGsiB
tJwdOc+CTCl5Egjxp/vJQXvTktbo9IFC3d7a7pu/yYw4/8J7/5JB8G3CCHtwU5yF
qnh1fGI3vqmDyzgOd1cWXbNVI+XN1dD/lnyzuVhYqHT7jfF2zN06oexClmVLTPfC
9LYcojylETJc1Ct5KpMza5w0ysHyZl+Y2Hp5caSrc7RU9OUb6opSF/jdy3MncoSO
weDGmKqpzLlAYt5omY9GEAdT6INsMvkon1gQ2gTDdPxzI44gMNVbcN7yW1aUG/nT
URb5Z/dIzQ+nrHmnywDVqDUb0ucKschz2FAmupIeHdZTXwYbJblwLZKUBWdQ7CRU
Sxrq4SGqJ+zG0EVw05IPGU9FmUF0aeDuyFHyv4Y8hOV3VUADnD0b/Pps03lgwrOJ
8vQOzGDXigKmvNAoejSIwEWmLuqbuYi3rKSZ+SKetEkaFLB5m0TWQPrI73OHlNCB
lbA/iXkMzw7bMogfI02MKU6Fw9VHPJwLUHXLxV2niQOgYztQ88aXUZHCt4Ds8rtG
ubC0iaGy9vCqfOr1+B4v/INyeT3fk7xbn+/MIBldKxr2ybAD57w8y0DgoQQSNssu
fyzH06e9D4OpPFxny+32z+rUku5s/SfXOdCIq3Nb+C5+RU8TdZi0hNN6hQuo0ylL
4aZBrzJtX9+/4rklzfgccOT0BIv7FBs9+9dQIzu6MmW2/ioldU9pM7a4RutjX04u
OFV/J4cfQKVKYo6ASxSpVMtbNVo4JY5JynP6RluUEtl6A5hzEheOiDYRZ3mxEFI4
01zU2+80XXBkc1k4Z2qoCyC6Hhoj9GuItbaxZhmbVsDBP1whM14J48b/PMbPjpZ5
u5k1nSyK2VVTKYPyBEf7GF0MlZNWeFLmFAVIJJqaizGV5RGeSxZtIx8jurx+Eb0o
mkDR9itR18W+BzcQVI7beOamijJxd4aaPKMosLuLPNFd+0pXth26RyufPlbaiRLu
wIHrJfyDPEMItLUh7FyGJpRV4ljGY8vmLThMUrA9H0mWnAy9VLYC4Lauw/uEg6CQ
cPgclsmIFtdWFF8JxBeOwrKM2u+TnCkrqiomgxMbADPYBW1Z+3O6GrWi827/5Tny
IKzVJGsEo3RmCu8FDMZU/mscgE6xGRrWbKt/31fcH8s+BLdvBtTGhlScc+zQVcGZ
bTOXbcWMtPv7qXI6AdnOQeUJ5azzIuDSZrQQiRbJHz2EWKaA5OcyZXHuEObh9ay5
3CFCI+t8sxy7gKswUmDG7PvcIcs0deUaBXSeTxEl9HmU7Rt3LKJTXvPw7J/Fhc84
a7hsPn651cKUQ1VDqgnAk8OGDmlWpf0dQu8Gl6XVB6OS6UeOCIeXOA67tYp3yx/A
qCE/WrPhCBbb5Z2aE75eKjMMvxtDNXVGNqyGxpnpXoRUJ6u4Mo8yitgqALap70EF
koX9Rl6I4lwlChOGgkq8QgIJK/C91PypQx/P/miRs6GCESDM/QGNyloNTc1Dpon8
3fArEtJP6EaC8ZexqIKbWPuHcJ2Z3Z3MsaXJWGfwbsCHPS5EPBc94ufo3/VWGld8
Sj1f9ux+2XB42Hg5sNBgBh2xnX/l9dpx1+yBb4nr7ZLB3XC/TZYf5m1MLvcnGqGc
v3JVyDejpjE3UfQP1DMcTIWjgAXcyV7hgKOhm74Lm4JhbKwM6lidY4D3lkTG4T9o
W5gQ1kNY3MtlDRhx93IWmHrrwSrYtHsFhY8dTlhKeRh73Wgxh6Nk8r6qzOi1EZ+v
bKGA/HNkuUMe83PCwOSwqWDnBKNbwhhaSn0yoKDkJA+vi8VeMzTBKHaWchoygqQR
iqPQa8sFFGrfRfo0HBgGiIP6/9ze1fbaNRgbLn9MUlhvLAnfWhUEb7dU5aJ9fWBS
sYHuNLg5WxfrB69NRbI0VUsj+G+YStN0RCzaDZz3az4lU8ICWBerQ0Jh8xBQCRhM
GglNJKbdPBS4wcyYydy/VfFANZkDH6K/X/XPm8CfN3uYXJR69e/OW1qAbJjtYVuf
BSJEjKSgjB1lS8NWMBplkulEhR07iHH9JEbht7vZ561SScxAOc+MmfEiP4qTEFwO
TDBXiABgIrddq2gqE6PUJ83ITNS2pfuS8hgvtHpzPLbwxP3fK49nTF9F9V+qhp82
nR2jbRYHdz1d5uY4zrQuArTbALRz2WfgQRfs0nD+MaT9sWavfxhUsbre6dt7ZEuG
bbNJNL1aTvuJv4VJHTmpM8vFBUjY2Km4BLpNOfBJe8H/574JQtj1I8ETS/YGSLMC
mPqf0N2Wzvxj8sje3Pnij1vry6hfwpuMkXdBPGqOwUIxHvUL7+okBJfRPIsyrIOF
lhFQFh2uycJ/5M9jOgsdic9zFQYBzp3DexwPehkCZQUGBfMylxp2i3G7KbT+JqJd
Q08Mujqaoi5WoMdmYsZE/qMmyvGis7C5hSsmq/6NeL2ACXY2VvI013JhmtrTdryg
SwHmFirwF3QcS0tGj3TQu+LrEDqsrve+6opTxFvwVMuaumuKM9vZrkRT55t9E+EQ
DhZbis/PGmt4w1D4KfxHCDKCxzFTH7nkVbPVLnEVDjFk8sH26vQ4UMb0abMnEi1S
JJNN7XFJFv1vHDZYIwl9TDws3V3LiexqpWCRLRVhJ1MDlYv58H+BF4VvHxZrsUmd
/Cm5SHfOIfTRypq7isZcOJFSL+4GOerMCPUcKKHo7sIesmdA+ePfpbkA1IEJWuRX
zIreJxC8jCazVPG23edz09NNLs04InRoCPB+F+L3uZh6WQj7RUtyCoKTlxkRNvXI
U97y3HtJgJ9aZBXyXa/SZ+rWnAy6XEZRb3PZ09H7ObpfvGnfZu159WK3QN5oM/wl
DinAXHhu6ZxOfZX4GxnHVjQub2ZgaR9t/1vQFc0fajauTHvnjiRg62d+D+UmzJIZ
wI7lZ8DMRcSqHGe1cZteR29s0lGXgpk28tIxnYnSyl+MPT7nFdqEbFSztykUBzAX
H6gIf81LpbM+qGKenIA1u+iOnp2fG7hB7OlsX2ZFuYh2HAqAnqy/XTy+ZcGLZJ5O
mwWyDH5u24VraCQ7t882YKenxcPmcf0IDc0ogPU3lQrIpDQcHQlPCfV9v0M1ulGO
OEnfZKlvt9m4V0BaO5dWSDcODO1meaOXuIh0k5cSHXawaUN0AtKc36yiv6gN+Wim
SgmpYg0muTtPKjco+gZNkPOq7XflLGxpzCiljJG7i/NUxjXFgJ/onZLOqA7fsE2R
k81/PLhYfoAdEcvAPjRPm96ExW0+0YJdfobJ3yJ5fCindIDmD8saFNUJ+dHzXl1h
eCDdVrQuNeUoKHyrqAbztw2Ju4zM7mSMhKPOIblhZVliqYP3cVsVaXwTrBULpK5E
xc3jXHZcgUPfyijxljU8jkUs5Vyh2CwmaU04HODLF2KV0WlXoovzZ6TR68w3O0bV
s5aA1TyeosNf4Thb4EJThDS9kKqyrAUUciEXEbkb8Jewd5EDsNT2Xr4hGzaXTQc2
lUAgptGxB4mBm9Av2NoTmMRCOGls+EBD1WFC1lad7Bpgk/utsfh24OqaB3LTONqZ
zNT5bDhmdcU2r/oI85M3MlvAaDFB0x8ZaZ/NcqQJrPx98LWPi87OTq2AjX7gcXtf
msTvRvkeWNd+7i26TeQuBD/ad/HqQsTW9IJKvDqd73abImrhdS/e213DucXfLx9L
9UYsh+y0GtqVHtHqlIFrHG6HPXgswrRhAtLaRB2kv/64VHVBxStTgz0a29pbhA4+
ZOCcrZVQe//osN5jcCeMpIrcmWh7pqUOTPmUYM5LZmUESXktLU+YTQAq9YL4copI
vRrNfasD4Zvf1HiIMUrpufp4TV9UIf49IqRFhk52eUv6rfQ+shZ9cCTAdT77hw8N
FeEiRPgkrzIUJPh8wxwi4wEhdzYAJnAEZTInqOAXxAYVVJSxXwMP2E9GBlEglYbi
77VLTYAstXnZyHhT0TXwe/d/g5eCFs8Lm2tUAv/97FEdPeSRnPDobH1jt+90hEj/
aGmAxLQo/cVlDOmIuoJM/C0Y0uiWfGV2gA2e8iEo7dD8pSKZE66PwlFIHi5/C6hW
BNcJpu8a6WdxKQRDqPOPcXrmYv6Ki0YUvxJJ8JOBbszpcAupOStMR04Q/9tuFZah
d3NiYTUjuBMFGUo3WQ5K8j7Vcn+zUCUxM+3PoYMmI4fqiJ1/3fdSGUYj/EGiBorr
4EJpO0CKPLl115YE44r8tDhiQjVPhb6A0G9ki3msbxYYI67YEPdZhBW6HNauYA7v
Ou7kPQ4yhXFNPXfff2Kty5tUmtYMkm0PGXv2roA+loUfae5ZY6Vvor3Nf0wjkSdp
38NfPlE2ZY37s/ZETI7sRjfq7VO7mLXw28+7ZBrqCOmQCv7Yz32NkQkQccaJvxxr
MXdY5qN9wPawV31IDztqTifIA2HmMrDhdbxkSv62NQNRdcIUXDA2Xb6aX6ro8vM0
Fm081aBslawB8wF6VJOGIMKNaSU8s9r+Ko8cLvxv+p3u/FEQPPaA12ysos3VIgll
/x89HccrN/aL8k2B3TSKmoYzGdE6b2t5hZ36FMCt3g2fErlIq4JDz0b91KU08eoU
5bdMXIGgeGt3wHTNcnWjnkXM6rCus2E/zT0LIjSdpn7qNxfSM87nJ0RdUfXcOIaY
9c/t77/JyMj8ccvSeDJfkg9szkN8oYcLUeNjB5qv/mxm5pJqFSrfgazw6l2/X3fR
f88kxo67ntlTSJFeevn7UQ6YsL3BHhokTupYJKGLj/Ni/ywtOiIEqhoC5sRgqABr
eur6NkQ6me0fgRDsR1JPIQ0aWEPip4I1NEBZekcMjVlxRvqqK65I4STuM3mJtEvN
Nm0WDKMx/9A+8Sx7jSdwLiDTz3ewzvSNy/Cp7dPOlVLhFMFBdfzkttRQBAz2aHwk
4iHJ721sdOkEFtaJbP4Mu+Xe/2QWNMbuU01YXMiofmd3dBYX4cAJUSRSXFReKTkj
c7YHT+5CmK68NjBzbUd6I7elRvNLFxURershZGLzEplQfYxgfJZ8B3p8gA+xqHzg
oYSVb9pXoXtkQeXkhI7J9e9+tvKKgytLXhk9I3zDEVYnnZgbLWL9uWvxQIMWqZoZ
vr552GJy4ybirNaR+s5biJAiVbcOLBuNS/Dqp9OzTDToCYm7KLP1AC9YHHH9V0YC
+b5WqdhtTL37tnLJ9VtkEToedElLcNnr3dySm8AmyAZwNL6+qSoiLfLlVoZM+lU0
cxcjkqG+NFXrT263IXHmWlg7hsEBiwd/xZIGUMsNxjnXQigHBTOyfBO4aPfrtmY7
e5GQ7CL46hPoGGRwvoTSEgiqdQZt2a/6z7tYSNxU5f32AnPl2Rb+/0/+e/d+oj64
Dv2BkxlPlfq4PU1ImQZe8zzH38VEtAymoSc6LmsyPRUEtGJqQXUlHva54q7tWcYl
WsugWu3BIWroDZUuu6RNxfzORU0xoNGx3o3CmN9PibNUGeavnLnBMUVtNhJ8LvEL
aASp1OXTPG2CBRxgnfz0sfdLsVkjqC1bXoVKEn2L9fKiqioU4HOq+OmqPXpReSxK
kE+zx63bzjhrW1Qn+GQoGCL/gpZSZVjBXMnhRDr4zZBFw9QtGjq+0ikbBjDtU8QS
R+p7TjYefNE6Hc1gZ3pWNTqa5AePcCkS2Bvmt6heXsV5+t8PTly6FcAKMOmjIHdF
E4CPTYdh8LwdfvvLy8z8J1SY3Qz6DHozB9FIBXAzg0xs2keLCG1+XTEIyn2bFNOT
uZlFj07PYEoSceJo0az92DQk35uYAHbciqre/CDSS0pf3C/L+LQrGoAejQIxJ3ff
fIc/v8U7TZ0s0Ngey/VW5n110fWA5ZQzkziiq84JWx23XNiaZ+vrofRY/P2hhWdl
XYEUMrSHfECwD1Cu45pmZryPczwFLO9pm64DM1nhjlV26qnk7VT1u22qhrhsq6al
yYej8Ls7exok2X6K2sniZphSY1gZJslyQwULeQ55Y/nZQZN4eJ74hNgSeKGouEdW
fZyglfg0UVicnJhLw9gi/dxqSz1dKtAybjsufSb8OU5CzHu2lOyZsVUgVzL4fY+l
816YYv2YQmFxsvPoM7kkOOmfS7tJb1/aMoGXvniAFo/Ptz4EHMFSHYAJuQ4DbgK0
6HLKI8bWDavuXHnX86vbPn1sOHhpjOR/psF2+zLoRykfpEA7Xozedp/jnuJoD7W2
UBtmDFF1eYPlHinDSWhOkBLLwkU3QUSlpBVy/+yx2dFZBGv3lrhyKAwG481L3liE
wVEi39fu2d3QDFBJ28xMzdTQ07kX1F+xCluldreAYknBpRn09sZJMBxkLROGugSy
m6ad3SYzmmzbhkYqMhx4a2q1JUkZts4XXBo+S+SzgHR4Pp0Lt7TbeHqUU6AGMaNr
zf5kOtATUVrM+aWUe0XRR6XE7gRLKhBwOlQtdRJ+F0nW65gqN7y6YcqWTdmV861r
9c8NWTcqqjOirZNd7R67+Cb8iWaGfylaWFVn0O7LTid9ERQDCohlq7rLDbrNtA0t
tScxdMxcWmIijmDH3KwpaSfb/rm+R5/bS+5Quc0GdoDmZZWNFVckZ4RPboBnfpTp
S1zKXOV6WjGjwv7yNrEsLBms1o4YZ8dXfVUPStXoexYxVA2S6I4ZSG9b2QHnO2PN
WGfnAbJ2uPr2x3MHHxE9gHDAM+EhD3Jpou2yxtnaUmSUdbp83L2bv5Na/ntCurmO
RpO8F0yn+JrEivVOLzv6i8JxKv01vKVghSMD9+YOTTLPZNiiV/BL9PL+112ONXJR
MbuL6Kr8nkWUSo31n0/PfENUQC+c/55amaTOnm4Ex9eRziB9lA8lV4857iRJ0t+x
9XUwq5z7wwa2cbb6cUSHgmab+3JZCDMA66Dv1A62u/U4XFk/XXSRPG2E4VmPvWA3
uQPSjJ8KlzM7k6u9sdCeRE/aPL1A87CI6GBbwkss+J9hsm3ymDqdyKjwbJlflF42
CBuazhl5J1xGb+dSDRIyiQXjq+EpVKhNsxlV3O8rdqI8D/zCg6egWeqlju4T3SsV
M/QTowq/WMipYI9RUAU/ARkOkA4Gq9Pj6U4jWcefaDDAj9RlktdDJeEPLQ36HiL2
ui2Dcb+fhi3V9Hcz44M3tzKFhj+VmvYAXwndzN9u6Cbpqmb9RCfZSlFSN8bBEXsf
EaC6cJWXn5h1iemGdxlmPMGCzRJY7vE01egr4y2bPB2lPfLp65chw5URvZ2vn2vh
lg59BnUU9/D6u4kMZA5HFnjbRZj2Dc1r95SpsXSB+7nm1Xw21GVyAeyvcceaQX7j
pnEUIEzL5LhXj8w/sOma1/jpibqPSDOp93shzcJANNube7B53FHI4MvK44R05Xb1
cN1sBJ1ByeXqV//CFXoqRCK1fkrX0G8u/RnAhMusehthjpxZXuQOq1e+Dtw9JAwh
Hd2AWhQ0CbcoiUSCtypX7rYgdUrm0Gt/CZi+w6DWkO8SwpE+JS4XhDawoW8NirvP
rUDrkEqOz6hh6/c2+UqnDIZFGLt3kXSAV4YFDDb0DFELb0G+FnQTFwCr1WQG6yEY
VnIgiBvzuCwbh96XPRev54rDFQKMflGy5efQgsrf9uLPRCYpDmPIJMNAWpO0deBR
3PbSSbwPkZKeFkVfmIqyhn+yOtKx6EVyTu/4s03eYdRq15SJfYLbYcD7evBFD/fB
q5OiGzQdd7L8XmsFgAmy8uo7ovPlA1aP+yS5XuSugLTxTcp28a0MvkOcZj0FPYaT
VAIFJrtJRbXu72U8axW8pU8vLRqv06rsgAHvDbZxIACLVAkLejN/aI3fIRh90BlC
3DmqW473ghSXKW/RfVT7KKnvN1pu/QY/MIKWWU+L5OMB4n3dF3XeSDrK9gVbvO9U
ll9q9Lx/8O0qU3wQZ7+peWCysv1LQEKHeEf1fJvIl00HsstnDYcvSkseYpP+JBQB
fuWlpknskY9IGAd5MShE0twAnxNQmWS6pvSnV47nhV3RKr9W9V0xQ9sf6dqEn6lM
hKXhvyYxpoQcqGXqCtfM7aLwG3V35J0G714pS65v9Yt8UTIgKvdtHGqD05L2fvFq
UxoDWIWeYxyTpYJmDd1yLrX1NdmRaeP9uI2JHsCVm28paiiE59528ikZbr1x8AQb
Y/Fva9ZaAQAw8sgr3YDwn1EcQ0ZWTrnpfkTuxaQLOXvlgInERwc5dk6AOPoIAw8R
Y0EoiAMBIfq/E7/vFeO1e02XGgjKsHU0Dcr+cmpMkY3tbpaqr9VY+hcGUbUbgwHw
Y7wWIv1Xo2QRpduDyNeytLgPRjvKCvz0SDuBPDeh+WwtmeFw/Z9E/qOj+0gTiJ4o
6EbcRQnRWwKiBAsydx/sXs6F0yVzhBl+YNLmEKILiV3M0PgruY8jMbS+1nS8GosW
ocGTCKNNMI/gGrMXdXbFl0zxojOgJy84AvQd+y/zFw1UNTRRNbq/9YvadzcUgnGk
v+yrFjCc5ip0lS6lcrF5mJ8xLLzTOWcA3IASHZw37HD1Qx6ywn6pqGijigVp+oUQ
ZGtGiGmYg/K0dpqrn/dhgnWOHcW6F6UGcrruK1Xh/B7c0bHqbrZKIozY53X8sRvL
VhghGzymJ3AcTJ804jvzBMwo5al/uytNhtvTsOw/JLO+EC4BzC2KP11ooUV9ajoC
bPSrODcRmZsM9RjW7jyF/gVWKwj2QolWGGFzef0ceW5WamLovFehtygCjjZBN3OD
YLJ+l4V/HeUwUuD1itNvdnND1Hz8RpGeolEIUbQMN4dfjitwtWG4cm7OqggMwUBR
REcHKnULY46dvPF3/RvVQVVudP22D6aO5bj/bVY2UZsr5zQA05wI7e5U42CZiI23
eEQ/nvAdpCzb/0gJLkfjFtuXvwUgIH/hwfRUzfGR+bxyJbapWS6MfwEoOr6mK7VX
0Ut+QBoPT+snliQQT0gnVBYgAr1JLHJyQoXgxu01xvCVJH3LQdPLIweEPKTtQz9y
MOh6/D4PMdMSkmzYebf4KeB61Bck3FuXYpfWv6OlYzb6Tn9dozrk1sDcmg+3ofZC
FLe4Obw9AwPLWSsO4sMmjCXuLOwYw4DdEXEiso4p8k8SFuizpF9TIANQPKBA9/MF
UCkZHXp7GLALobgBHykgOFrqrxoHza67fpgkAVcg6pGHlKsKQ1QNOLU2HHN/NyIx
lzKQf1yNSJ6Q4W4SvBYgLXUdHTsHtqXP3OtAL31RgkLO1noG/xDA1O+9khX2YfaU
yQM8vVk32A3fmx8CHKzrWR2wgGPujO6rfpqJ8Kpg8ZESDbNjpBecMD6SA+H5nLsl
JuTS5hXufOJebijctMquxA9PUhwe79LEUjet7rViDL2E98fx6KYUz7x73cmv3kIh
9dUU61WbicNfQjAj+/9hc6hvLOLuNJBdyiwDgzM/K+uv3kmSVGSPzDPUFSnmf55z
QCrvn5rrjKB32D9v6BocMfeseT5uNlwDsI5//lXGvVJUPgPP874qKJi9/DYyXnAN
fKv4bhBtyZjR+wkhULtm3KWpFrWqzpeG2FbowwC5o0HPCInB5WIBW+Wozi5guqOc
PHViyKonFXgS0RFers/HtAN0nrlWTgHR2oXK7EXUNbhFlQgaTTWgtuUzfwSWD+sA
oDDlsjj2foRmfAVLzHAKcTrGqlDtwzprPJfN2fJbFVZLFxDcDUsQwNzFVG43H60z
IVZy7WDw6qfhHSfYTHiBIFaYtUPoWzY3yS5Bi6/Q4qLTlG+/6Y4/jlqpav/TX4z0
lLjjVzDG9X8jnaWr9wTiSHWwpCZihr2FjFK3IpTQhFo8Z17m+7GdIEiu6GaPo3DD
FPwA2kqV1EE64NUt0geCO/x0GXrEQMnf8SrkaVdOtiWnVOwhAfK7abj9+18gKj00
2qL+MaeXft6yzDYPkXEhUDdeM/lAIYVuy3RiAPx3pkOf9aniqUYe/+VzzCMqBMNz
S9GW3v5DSBtvkrRQF7Fai+TVdPeN5dZbKy59pJNrZLCuZCrjVXMk7smMcBPMv1Fp
y5jFi6DYfcTEN28dDbmeLgcfj+64s9PUiJDjGi+2GM5IzgRvKtyL1DguZTW9e06X
V6rM2qUXFjJiNxeQ/dCYFUnPOdCpUDBQyHEy2D9DdlINVuBotgTc3z6oaTBDeKl5
mvEa3XF6jVas6rasftqXZckBjzDC9cQv1pJcLDNLi0EzUkVzvJDctvIBW05ljig+
yLU8zDHxDD/HeNSH9/cHu2HlmLLHVC4I9Ek5XRgUP8IcIWt2KthsVcqkBi34Zplf
IyLFmeOXGlGs00529fTqKrH28gzUO4hSMwT0R312qrjNQ84a7dDozEMOISlzxk/q
Hn5BV0lcoK5DNCLDCbV4Nhjh+vk8bVnK9STKl880ZgxMo8QSU5pW0R/2oxN4VfaH
P8x3PqPDbKqqlUrmtrXlaonnTBlT3ezgaKF1jIPLApqxhTi27hcPj1SGJqeb2sqc
FZ+orqC1MncUO+aly+A/MfjoofXlEKTx9r0KNz8DXGD7YixB69S3buPo1S1JS/0D
MCR7S2dDftXTyrJsY77lr4a3J3Y0+2nQHA8md+tv7Ma6Xy/EG+73mn++yk1ONBjY
SMsQm3ipSrFd7LvlIbG5YhJy21kBPh486Rgl1ZPH/+86l6VCWxX0qYlGfypmNi5/
A8rOUSvEAty6wH+xz1ifCjeUG82Vipx4NZe5DGc0+uYQtunyNJwrfxaNxqCPLNUh
KDQdU5Yh+zISv+6Vj7mKf/YWOGU5ZGJ2cUgao17vx/pzNUBqLyqt1iCfLp9ewWsg
X8NoEpgF47XhvwXHS0OavyyF6iwaeIKAqWGJWQG64rPPfiiuiGDZefQb78cpIZbX
SJmSGiSSqjrPfMwPu2/wRq3pTIXv/3bpnldYhIwIW4FvUSXDlqGSKOw5Q0Lz9X6l
XOBxkbBboiI+Bww8DXr1tSCKMOc9qwy5OAJm3NS6XLPqGY2b/VmokwRCZfbv0hhh
qA3E/qL5FaXOcQPWsIIlmtrnX6JdPdfYM2VMC1SK8gKqrp9uw4uViLV68l5y4e/n
iWly+8G25SXLtgtnDhTYoPY8aoHmkJ4uasggVQZgyyMB968tcTW8akjnCFGdhySy
Le2e5k1wn7BL3yBBEkCEQhTiuF9cHOa1h3haepsnGTXeOx8LCbnwkmXh/40QBgx0
9EXjZi7tlpDHpLSRTUr/ftsRLIKyELhMEMtbbJgvN3308n7kbDMmrZX8GY5ZC3uq
IX9Wk/yfpMcFEbpfTyNSvcPElDH0CFS+MQaYEYPaoeN/Y20aS1XqNqX8npG1dP4G
LtfDfr4ASk8/O6xk4lmnAestrl+bEpMeAv9wOYPdbWcqFXgmbsI4boUsAp/LI225
Lh+BrFUcWpPUU2Rum4kYxCBQ6oKUl0U09tOcO83o7B7ACpyaIU1rh8YRC9Yl+1BR
jqf6yJm073bT1H5BzuoITtf1j6Be+CAQnKY22HCJ+eUeWLgX/HhPGqdoOT+uDwV9
bW/wWpqNmoVoYR9yJQJzmM5fbHxx/GeCLTup7MTCw0yxPO7b3/TED7rE934vkw2d
LdwhlCb4exQ79TB8f0EnYyuKYLAipE01M4L0Jj6ADbwG9pK169zRvZ9mB6oYL1wn
b/hp66YVcV0wbe77q1hZ0PRAO9FMsoYnyXDWiYO7SlOzwS8KVU475qnnHkN8ibEV
3anopOfdu9o0/a667bJ/P4vAiuh2o1Xp2cD7lH4YrQlm0MX2fHsbNCsi/jRTd8+Z
oIUtVJIvt9AFhulvYFEFFmXaJBBiqwcK4RpeYRsYAPKiNdplyrwRhcZFfzVautTB
LfgcqbZ4GKkD46Plw8iD5VoWEiEqvfWuSBZlzgjO4nMh07taLG9WbUPG0RBmlG/Z
JmE32D6VltVU13PMKMFYzD1dRW5lU2nFI3uRbnS+l8aeMABW2piidAkuiCmOhDtA
sfYEEk86zDKTjw3byyieyvtzBcU7b2L4DV8WJjAvwS7xnGFlfVCoUmKeQhvvL0uK
XEkTrMCOFH8woqDY19ABngq2pWuODRq3ak7Tw1gNfjZy6ej17sFd7OXxB3n1Cito
DSRnP/YCzSvQnjcVJTXUNpI7/eG9ox1msT/K/RT4CrSDCuFzO7kNcoD0tBjjkv5U
urGGJZlO4mZS+dEWlhOOjDkXNRTdCMX49LRXA0GMuRf0C3A9CKTke/aefscwNKxZ
56GzlA2EcxpE+Ht2A+fVpWlCxHrU8OTS55400Y9MSrVsOZy0NWLVmOdm2IZ6/bQ4
k7skAWyBObhk5NsjdODmTUq4sCF4KEcx2DS7MmNtvSMt1bfFJ+UoMDrI+XtIygvS
Nckvms3pzUkm0Ytvsf1S2XcSojzUtlaYgA3PT7u7DEmPiBLCrCe3X728t/rEqP5R
jyjqn4hXYwZbHQ61SZD9Xam+lO/eBNl8y2VdTSaki3Ob9E1sdGFgYia+Ek2Atc8v
mnJwAU/I0r0Ie422BP70Mf8d8maxUz3uQrOGUkxjEIctIo33Z8z0MdWrsg3edftX
Og7ukaAHeqalU/CRpShYxHnK87Zd1rZ2qtzu+p/aB58K3Ykzlp8Bo5gJYboM7M3Z
GswbyTu1ZnrcnvJogiXm/jEa5/vqCUEoy2FNCfKPNwJhPKRv7QaK/yU+Vv/etocT
SjzU3KzMd+g9g1QcpdAI/oTlTU4F2EFqJ9jgFxVpPDlRmXJpck/l49lsSX7GGAS4
AlkiCuinxx1ZdR9BfQ3I2G37h+ifLv1ozTyxHMqWdzyoK6C+cF6LuyCcpS0exQg4
c7A8tbtJIEmTCe83OxiLxbtu4cg7BULJn/bcNp5qeXeyxzvi3EO8lBpxsXNXHwoB
5p4VHk5tmZoornDuJ+BZ6bbV0RSInT0o5vpIB77SU0lAjBYZXLibNN6f0gd4cp0P
27ieN+XnarRXaPBb3uojWlaCwf88IH1s/L7e8Vf9+IR5H2fJg27Sp+Z1fHjaJi7p
Sb6pBXgEN0TJlEXpp6fs7x4dyorsakFWr7mHw7RWddJrls9fmcNQgjPF/TCvoiyS
RFbd+xvLoPoobS5PLbJ+J6YboR1zNlACmanHi5yjc1ww93SRYOSG/Jfg8XCnxOo1
oQenolRIINNyyS+FKsZNEzrddbJGJWddiTXYuVgqkBkkNrK6QWcSbU9OW54euSp/
LO4PKn0iIMnpvSXaXd4+6pBQMWZXEBvKXY8FKhvUNQJf1XkvU1E/JM4gA0wunxSM
yX+0T0a1CgGrEnDtK//yBwv91RlVz+K/U2JURVKzxQ+heGbRAGIecbK0mhIt+pZR
rXjaXH35vgucm49kkSrFns2OWFnMXzBitcV5paQbJR+P7jyywaWXvFqYKGaenTS7
QsIcdhQeajc9zDCmJi1pZK9zZrIeB2EXR/HUERxqp3A+1XE+CHbGhcvIhkVNk+t2
6hZVVgb52FMrfw9TW+AKekQZMkNKHVho4Ni7JzmujnU/XPsR/y32II7mcl316iex
hy9p61ah5An3MCvYi990vyPeB8ACWHvlYugyvmTYDJ61HAmlyfRpZpEQR0V3qzfA
s4+nV+5rDHqwnEo2QOMEO6qg4lJH6n/TfcXh2M3CBKSyzLUArlj1EMco0iCFv1yn
o+tHp92kfm1n516jFumA2yEgN/p7txm33Kt1GGivvfSiWxD2AdGV5rDvR7IHACU2
8t2GxNL3OCU+ltfjz0ZehZmt+VDicZMvPyEd75+dtCmRo+QHF4pnSI4+EJPCp7/p
CUmqBwRFGZvfPStbYdZXgonFKaEWY22XFW3pXQb1jMyu443vwmaVhYCErWSbSdEe
MKg3hoMLQwb/wiHajN1yfWsLUXR/MHO+VKIWl8Twoz8y3J87yu94EFFtwxqkqihq
aAnLwy057/ywOEkrCpCXYpI/epMa59sQAC+MU1sLvhZBiw66TM4SlBFKLNlrhOaO
cCjk+Ryfwf4dnozCkZj476TrDDgaBF5GeFsJJGYCrPFr7AYHKhL5Q6p70J84qN0r
66XdA6QWVo7VsKM0xApwPPrgRT0uwbny5DlT+LDO1xK514Wtd0s+eBIOWWNvJlze
gRSb04xPLRfd/e3dtccVcdXfyNn8cBcKYxt6/wC8qMSIJajDt3AVt1vVHvIQTqGS
0eM/kv3F3DaRJcqI4Jub+w==
//pragma protect end_data_block
//pragma protect digest_block
fNOiAIgRZRisII0Nb+YVv8DcspQ=
//pragma protect end_digest_block
//pragma protect end_protected
