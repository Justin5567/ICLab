`include "Usertype_PKG.sv"

program automatic PATTERN_pokemon(input clk, INF.PATTERN_pokemon inf);
import usertype::*;


endprogram